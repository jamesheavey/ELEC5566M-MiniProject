module flap_1_neg45_rom
	(
		input wire clk,
		input wire [3:0] row,
		input wire [4:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [3:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		9'b000000000: colour_data = 24'b111111110000000010010110;
		9'b000000001: colour_data = 24'b111111110000000010010110;
		9'b000000010: colour_data = 24'b111111110000000010010110;
		9'b000000011: colour_data = 24'b111111110000000010010110;
		9'b000000100: colour_data = 24'b111111110000000010010110;
		9'b000000101: colour_data = 24'b111111110000000010010110;
		9'b000000110: colour_data = 24'b010100110011100001000110;
		9'b000000111: colour_data = 24'b010100110011100001000110;
		9'b000001000: colour_data = 24'b010100110011100001000110;
		9'b000001001: colour_data = 24'b010100110011100001000110;
		9'b000001010: colour_data = 24'b010100110011100001000110;
		9'b000001011: colour_data = 24'b111111110000000010010110;
		9'b000001100: colour_data = 24'b111111110000000010010110;
		9'b000001101: colour_data = 24'b111111110000000010010110;
		9'b000001110: colour_data = 24'b111111110000000010010110;
		9'b000001111: colour_data = 24'b111111110000000010010110;
		9'b000010000: colour_data = 24'b111111110000000010010110;
		9'b000010001: colour_data = 24'b111111110000000010010110;

		9'b000100000: colour_data = 24'b111111110000000010010110;
		9'b000100001: colour_data = 24'b111111110000000010010110;
		9'b000100010: colour_data = 24'b111111110000000010010110;
		9'b000100011: colour_data = 24'b111111110000000010010110;
		9'b000100100: colour_data = 24'b111111110000000010010110;
		9'b000100101: colour_data = 24'b010100110011100001000110;
		9'b000100110: colour_data = 24'b010100110011100001000110;
		9'b000100111: colour_data = 24'b111010111111110011011101;
		9'b000101000: colour_data = 24'b111010111111110011011101;
		9'b000101001: colour_data = 24'b111010111111110011011101;
		9'b000101010: colour_data = 24'b111010111111110011011101;
		9'b000101011: colour_data = 24'b010100110011100001000110;
		9'b000101100: colour_data = 24'b010100110011100001000110;
		9'b000101101: colour_data = 24'b111111110000000010010110;
		9'b000101110: colour_data = 24'b010100110011100001000110;
		9'b000101111: colour_data = 24'b111111110000000010010110;
		9'b000110000: colour_data = 24'b111111110000000010010110;
		9'b000110001: colour_data = 24'b111111110000000010010110;

		9'b001000000: colour_data = 24'b111111110000000010010110;
		9'b001000001: colour_data = 24'b111111110000000010010110;
		9'b001000010: colour_data = 24'b111111110000000010010110;
		9'b001000011: colour_data = 24'b111111110000000010010110;
		9'b001000100: colour_data = 24'b010100110011100001000110;
		9'b001000101: colour_data = 24'b010100110011100001000110;
		9'b001000110: colour_data = 24'b010100110011100001000110;
		9'b001000111: colour_data = 24'b111010111111110011011101;
		9'b001001000: colour_data = 24'b111010111111110011011101;
		9'b001001001: colour_data = 24'b010100110011100001000110;
		9'b001001010: colour_data = 24'b010100110011100001000110;
		9'b001001011: colour_data = 24'b111010111111110011011101;
		9'b001001100: colour_data = 24'b010100110011100001000110;
		9'b001001101: colour_data = 24'b010100110011100001000110;
		9'b001001110: colour_data = 24'b111010110101000001000000;
		9'b001001111: colour_data = 24'b010100110011100001000110;
		9'b001010000: colour_data = 24'b111111110000000010010110;
		9'b001010001: colour_data = 24'b111111110000000010010110;

		9'b001100000: colour_data = 24'b111111110000000010010110;
		9'b001100001: colour_data = 24'b111111110000000010010110;
		9'b001100010: colour_data = 24'b111111110000000010010110;
		9'b001100011: colour_data = 24'b010100110011100001000110;
		9'b001100100: colour_data = 24'b010100110011100001000110;
		9'b001100101: colour_data = 24'b110111011110001010110001;
		9'b001100110: colour_data = 24'b010100110011100001000110;
		9'b001100111: colour_data = 24'b111010111111110011011101;
		9'b001101000: colour_data = 24'b111010111111110011011101;
		9'b001101001: colour_data = 24'b111010111111110011011101;
		9'b001101010: colour_data = 24'b111010111111110011011101;
		9'b001101011: colour_data = 24'b111010111111110011011101;
		9'b001101100: colour_data = 24'b010100110011100001000110;
		9'b001101101: colour_data = 24'b111010110101000001000000;
		9'b001101110: colour_data = 24'b111010110101000001000000;
		9'b001101111: colour_data = 24'b010100110011100001000110;
		9'b001110000: colour_data = 24'b111111110000000010010110;
		9'b001110001: colour_data = 24'b111111110000000010010110;

		9'b010000000: colour_data = 24'b111111110000000010010110;
		9'b010000001: colour_data = 24'b111111110000000010010110;
		9'b010000010: colour_data = 24'b111111110000000010010110;
		9'b010000011: colour_data = 24'b010100110011100001000110;
		9'b010000100: colour_data = 24'b110111011110001010110001;
		9'b010000101: colour_data = 24'b110101001011111100100111;
		9'b010000110: colour_data = 24'b010100110011100001000110;
		9'b010000111: colour_data = 24'b110010001100000011000000;
		9'b010001000: colour_data = 24'b110010001100000011000000;
		9'b010001001: colour_data = 24'b111010111111110011011101;
		9'b010001010: colour_data = 24'b111010111111110011011101;
		9'b010001011: colour_data = 24'b010100110011100001000110;
		9'b010001100: colour_data = 24'b111010110101000001000000;
		9'b010001101: colour_data = 24'b111010110101000001000000;
		9'b010001110: colour_data = 24'b010100110011100001000110;
		9'b010001111: colour_data = 24'b010100110011100001000110;
		9'b010010000: colour_data = 24'b111111110000000010010110;
		9'b010010001: colour_data = 24'b111111110000000010010110;

		9'b010100000: colour_data = 24'b111111110000000010010110;
		9'b010100001: colour_data = 24'b111111110000000010010110;
		9'b010100010: colour_data = 24'b111111110000000010010110;
		9'b010100011: colour_data = 24'b010100110011100001000110;
		9'b010100100: colour_data = 24'b110111011110001010110001;
		9'b010100101: colour_data = 24'b110101001011111100100111;
		9'b010100110: colour_data = 24'b110101001011111100100111;
		9'b010100111: colour_data = 24'b010100110011100001000110;
		9'b010101000: colour_data = 24'b010100110011100001000110;
		9'b010101001: colour_data = 24'b010100110011100001000110;
		9'b010101010: colour_data = 24'b010100110011100001000110;
		9'b010101011: colour_data = 24'b111010110101000001000000;
		9'b010101100: colour_data = 24'b111010110101000001000000;
		9'b010101101: colour_data = 24'b010100110011100001000110;
		9'b010101110: colour_data = 24'b111010110101000001000000;
		9'b010101111: colour_data = 24'b010100110011100001000110;
		9'b010110000: colour_data = 24'b111111110000000010010110;
		9'b010110001: colour_data = 24'b111111110000000010010110;

		9'b011000000: colour_data = 24'b111111110000000010010110;
		9'b011000001: colour_data = 24'b111111110000000010010110;
		9'b011000010: colour_data = 24'b010100110011100001000110;
		9'b011000011: colour_data = 24'b110111011110001010110001;
		9'b011000100: colour_data = 24'b110101001011111100100111;
		9'b011000101: colour_data = 24'b110101001011111100100111;
		9'b011000110: colour_data = 24'b110101001011111100100111;
		9'b011000111: colour_data = 24'b110101001011111100100111;
		9'b011001000: colour_data = 24'b110101001011111100100111;
		9'b011001001: colour_data = 24'b110101001011111100100111;
		9'b011001010: colour_data = 24'b110101001011111100100111;
		9'b011001011: colour_data = 24'b111010110101000001000000;
		9'b011001100: colour_data = 24'b010100110011100001000110;
		9'b011001101: colour_data = 24'b111010110101000001000000;
		9'b011001110: colour_data = 24'b010100110011100001000110;
		9'b011001111: colour_data = 24'b010100110011100001000110;
		9'b011010000: colour_data = 24'b111111110000000010010110;
		9'b011010001: colour_data = 24'b111111110000000010010110;

		9'b011100000: colour_data = 24'b111111110000000010010110;
		9'b011100001: colour_data = 24'b111111110000000010010110;
		9'b011100010: colour_data = 24'b010100110011100001000110;
		9'b011100011: colour_data = 24'b010100110011100001000110;
		9'b011100100: colour_data = 24'b010100110011100001000110;
		9'b011100101: colour_data = 24'b010100110011100001000110;
		9'b011100110: colour_data = 24'b010100110011100001000110;
		9'b011100111: colour_data = 24'b110101001011111100100111;
		9'b011101000: colour_data = 24'b110101001011111100100111;
		9'b011101001: colour_data = 24'b110101001011111100100111;
		9'b011101010: colour_data = 24'b010100110011100001000110;
		9'b011101011: colour_data = 24'b111010110101000001000000;
		9'b011101100: colour_data = 24'b111010110101000001000000;
		9'b011101101: colour_data = 24'b010100110011100001000110;
		9'b011101110: colour_data = 24'b010100110011100001000110;
		9'b011101111: colour_data = 24'b111111110000000010010110;
		9'b011110000: colour_data = 24'b111111110000000010010110;
		9'b011110001: colour_data = 24'b111111110000000010010110;

		9'b100000000: colour_data = 24'b111111110000000010010110;
		9'b100000001: colour_data = 24'b111111110000000010010110;
		9'b100000010: colour_data = 24'b010100110011100001000110;
		9'b100000011: colour_data = 24'b010100110011100001000110;
		9'b100000100: colour_data = 24'b110111011110001010110001;
		9'b100000101: colour_data = 24'b110111011110001010110001;
		9'b100000110: colour_data = 24'b110111011110001010110001;
		9'b100000111: colour_data = 24'b010100110011100001000110;
		9'b100001000: colour_data = 24'b110101001011111100100111;
		9'b100001001: colour_data = 24'b110101001011111100100111;
		9'b100001010: colour_data = 24'b010100110011100001000110;
		9'b100001011: colour_data = 24'b010100110011100001000110;
		9'b100001100: colour_data = 24'b111000111000000100010111;
		9'b100001101: colour_data = 24'b010100110011100001000110;
		9'b100001110: colour_data = 24'b111111110000000010010110;
		9'b100001111: colour_data = 24'b111111110000000010010110;
		9'b100010000: colour_data = 24'b111111110000000010010110;
		9'b100010001: colour_data = 24'b111111110000000010010110;

		9'b100100000: colour_data = 24'b111111110000000010010110;
		9'b100100001: colour_data = 24'b111111110000000010010110;
		9'b100100010: colour_data = 24'b010100110011100001000110;
		9'b100100011: colour_data = 24'b110111011110001010110001;
		9'b100100100: colour_data = 24'b110111011110001010110001;
		9'b100100101: colour_data = 24'b110111011110001010110001;
		9'b100100110: colour_data = 24'b110111011110001010110001;
		9'b100100111: colour_data = 24'b010100110011100001000110;
		9'b100101000: colour_data = 24'b110101001011111100100111;
		9'b100101001: colour_data = 24'b111000111000000100010111;
		9'b100101010: colour_data = 24'b111000111000000100010111;
		9'b100101011: colour_data = 24'b111000111000000100010111;
		9'b100101100: colour_data = 24'b111000111000000100010111;
		9'b100101101: colour_data = 24'b010100110011100001000110;
		9'b100101110: colour_data = 24'b111111110000000010010110;
		9'b100101111: colour_data = 24'b111111110000000010010110;
		9'b100110000: colour_data = 24'b111111110000000010010110;
		9'b100110001: colour_data = 24'b111111110000000010010110;

		9'b101000000: colour_data = 24'b111111110000000010010110;
		9'b101000001: colour_data = 24'b010100110011100001000110;
		9'b101000010: colour_data = 24'b110111011110001010110001;
		9'b101000011: colour_data = 24'b110111011110001010110001;
		9'b101000100: colour_data = 24'b110111011110001010110001;
		9'b101000101: colour_data = 24'b110111011110001010110001;
		9'b101000110: colour_data = 24'b110101001011111100100111;
		9'b101000111: colour_data = 24'b010100110011100001000110;
		9'b101001000: colour_data = 24'b111000111000000100010111;
		9'b101001001: colour_data = 24'b111000111000000100010111;
		9'b101001010: colour_data = 24'b111000111000000100010111;
		9'b101001011: colour_data = 24'b111000111000000100010111;
		9'b101001100: colour_data = 24'b010100110011100001000110;
		9'b101001101: colour_data = 24'b111111110000000010010110;
		9'b101001110: colour_data = 24'b111111110000000010010110;
		9'b101001111: colour_data = 24'b111111110000000010010110;
		9'b101010000: colour_data = 24'b111111110000000010010110;
		9'b101010001: colour_data = 24'b111111110000000010010110;

		9'b101100000: colour_data = 24'b111111110000000010010110;
		9'b101100001: colour_data = 24'b010100110011100001000110;
		9'b101100010: colour_data = 24'b010100110011100001000110;
		9'b101100011: colour_data = 24'b110111011110001010110001;
		9'b101100100: colour_data = 24'b110111011110001010110001;
		9'b101100101: colour_data = 24'b110101001011111100100111;
		9'b101100110: colour_data = 24'b110101001011111100100111;
		9'b101100111: colour_data = 24'b010100110011100001000110;
		9'b101101000: colour_data = 24'b111000111000000100010111;
		9'b101101001: colour_data = 24'b111000111000000100010111;
		9'b101101010: colour_data = 24'b111000111000000100010111;
		9'b101101011: colour_data = 24'b010100110011100001000110;
		9'b101101100: colour_data = 24'b111111110000000010010110;
		9'b101101101: colour_data = 24'b111111110000000010010110;
		9'b101101110: colour_data = 24'b111111110000000010010110;
		9'b101101111: colour_data = 24'b111111110000000010010110;
		9'b101110000: colour_data = 24'b111111110000000010010110;
		9'b101110001: colour_data = 24'b111111110000000010010110;

		9'b110000000: colour_data = 24'b111111110000000010010110;
		9'b110000001: colour_data = 24'b111111110000000010010110;
		9'b110000010: colour_data = 24'b010100110011100001000110;
		9'b110000011: colour_data = 24'b010100110011100001000110;
		9'b110000100: colour_data = 24'b010100110011100001000110;
		9'b110000101: colour_data = 24'b010100110011100001000110;
		9'b110000110: colour_data = 24'b010100110011100001000110;
		9'b110000111: colour_data = 24'b111000111000000100010111;
		9'b110001000: colour_data = 24'b111000111000000100010111;
		9'b110001001: colour_data = 24'b010100110011100001000110;
		9'b110001010: colour_data = 24'b010100110011100001000110;
		9'b110001011: colour_data = 24'b111111110000000010010110;
		9'b110001100: colour_data = 24'b111111110000000010010110;
		9'b110001101: colour_data = 24'b111111110000000010010110;
		9'b110001110: colour_data = 24'b111111110000000010010110;
		9'b110001111: colour_data = 24'b111111110000000010010110;
		9'b110010000: colour_data = 24'b111111110000000010010110;
		9'b110010001: colour_data = 24'b111111110000000010010110;

		9'b110100000: colour_data = 24'b111111110000000010010110;
		9'b110100001: colour_data = 24'b111111110000000010010110;
		9'b110100010: colour_data = 24'b111111110000000010010110;
		9'b110100011: colour_data = 24'b111111110000000010010110;
		9'b110100100: colour_data = 24'b111111110000000010010110;
		9'b110100101: colour_data = 24'b111111110000000010010110;
		9'b110100110: colour_data = 24'b010100110011100001000110;
		9'b110100111: colour_data = 24'b010100110011100001000110;
		9'b110101000: colour_data = 24'b010100110011100001000110;
		9'b110101001: colour_data = 24'b111111110000000010010110;
		9'b110101010: colour_data = 24'b111111110000000010010110;
		9'b110101011: colour_data = 24'b111111110000000010010110;
		9'b110101100: colour_data = 24'b111111110000000010010110;
		9'b110101101: colour_data = 24'b111111110000000010010110;
		9'b110101110: colour_data = 24'b111111110000000010010110;
		9'b110101111: colour_data = 24'b111111110000000010010110;
		9'b110110000: colour_data = 24'b111111110000000010010110;
		9'b110110001: colour_data = 24'b111111110000000010010110;

		9'b111000000: colour_data = 24'b111111110000000010010110;
		9'b111000001: colour_data = 24'b111111110000000010010110;
		9'b111000010: colour_data = 24'b111111110000000010010110;
		9'b111000011: colour_data = 24'b111111110000000010010110;
		9'b111000100: colour_data = 24'b111111110000000010010110;
		9'b111000101: colour_data = 24'b111111110000000010010110;
		9'b111000110: colour_data = 24'b111111110000000010010110;
		9'b111000111: colour_data = 24'b111111110000000010010110;
		9'b111001000: colour_data = 24'b111111110000000010010110;
		9'b111001001: colour_data = 24'b111111110000000010010110;
		9'b111001010: colour_data = 24'b111111110000000010010110;
		9'b111001011: colour_data = 24'b111111110000000010010110;
		9'b111001100: colour_data = 24'b111111110000000010010110;
		9'b111001101: colour_data = 24'b111111110000000010010110;
		9'b111001110: colour_data = 24'b111111110000000010010110;
		9'b111001111: colour_data = 24'b111111110000000010010110;
		9'b111010000: colour_data = 24'b111111110000000010010110;
		9'b111010001: colour_data = 24'b111111110000000010010110;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule