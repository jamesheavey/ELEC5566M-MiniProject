module floor_rom
	(
		input wire clk,
		input wire [3:0] row,
		input wire [7:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [3:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: colour_data = 24'b010100110011100001000111;
		12'b000000000001: colour_data = 24'b010100110011100001000111;
		12'b000000000010: colour_data = 24'b010100110011100001000111;
		12'b000000000011: colour_data = 24'b010100110011100001000111;
		12'b000000000100: colour_data = 24'b010100110011100001000111;
		12'b000000000101: colour_data = 24'b010100110011100001000111;
		12'b000000000110: colour_data = 24'b010100110011100001000111;
		12'b000000000111: colour_data = 24'b010100110011100001000111;
		12'b000000001000: colour_data = 24'b010100110011100001000111;
		12'b000000001001: colour_data = 24'b010100110011100001000111;
		12'b000000001010: colour_data = 24'b010100110011100001000111;
		12'b000000001011: colour_data = 24'b010100110011100001000111;
		12'b000000001100: colour_data = 24'b010100110011100001000111;
		12'b000000001101: colour_data = 24'b010100110011100001000111;
		12'b000000001110: colour_data = 24'b010100110011100001000111;
		12'b000000001111: colour_data = 24'b010100110011100001000111;
		12'b000000010000: colour_data = 24'b010100110011100001000111;
		12'b000000010001: colour_data = 24'b010100110011100001000111;
		12'b000000010010: colour_data = 24'b010100110011100001000111;
		12'b000000010011: colour_data = 24'b010100110011100001000111;
		12'b000000010100: colour_data = 24'b010100110011100001000111;
		12'b000000010101: colour_data = 24'b010100110011100001000111;
		12'b000000010110: colour_data = 24'b010100110011100001000111;
		12'b000000010111: colour_data = 24'b010100110011100001000111;
		12'b000000011000: colour_data = 24'b010100110011100001000111;
		12'b000000011001: colour_data = 24'b010100110011100001000111;
		12'b000000011010: colour_data = 24'b010100110011100001000111;
		12'b000000011011: colour_data = 24'b010100110011100001000111;
		12'b000000011100: colour_data = 24'b010100110011100001000111;
		12'b000000011101: colour_data = 24'b010100110011100001000111;
		12'b000000011110: colour_data = 24'b010100110011100001000111;
		12'b000000011111: colour_data = 24'b010100110011100001000111;
		12'b000000100000: colour_data = 24'b010100110011100001000111;
		12'b000000100001: colour_data = 24'b010100110011100001000111;
		12'b000000100010: colour_data = 24'b010100110011100001000111;
		12'b000000100011: colour_data = 24'b010100110011100001000111;
		12'b000000100100: colour_data = 24'b010100110011100001000111;
		12'b000000100101: colour_data = 24'b010100110011100001000111;
		12'b000000100110: colour_data = 24'b010100110011100001000111;
		12'b000000100111: colour_data = 24'b010100110011100001000111;
		12'b000000101000: colour_data = 24'b010100110011100001000111;
		12'b000000101001: colour_data = 24'b010100110011100001000111;
		12'b000000101010: colour_data = 24'b010100110011100001000111;
		12'b000000101011: colour_data = 24'b010100110011100001000111;
		12'b000000101100: colour_data = 24'b010100110011100001000111;
		12'b000000101101: colour_data = 24'b010100110011100001000111;
		12'b000000101110: colour_data = 24'b010100110011100001000111;
		12'b000000101111: colour_data = 24'b010100110011100001000111;
		12'b000000110000: colour_data = 24'b010100110011100001000111;
		12'b000000110001: colour_data = 24'b010100110011100001000111;
		12'b000000110010: colour_data = 24'b010100110011100001000111;
		12'b000000110011: colour_data = 24'b010100110011100001000111;
		12'b000000110100: colour_data = 24'b010100110011100001000111;
		12'b000000110101: colour_data = 24'b010100110011100001000111;
		12'b000000110110: colour_data = 24'b010100110011100001000111;
		12'b000000110111: colour_data = 24'b010100110011100001000111;
		12'b000000111000: colour_data = 24'b010100110011100001000111;
		12'b000000111001: colour_data = 24'b010100110011100001000111;
		12'b000000111010: colour_data = 24'b010100110011100001000111;
		12'b000000111011: colour_data = 24'b010100110011100001000111;
		12'b000000111100: colour_data = 24'b010100110011100001000111;
		12'b000000111101: colour_data = 24'b010100110011100001000111;
		12'b000000111110: colour_data = 24'b010100110011100001000111;
		12'b000000111111: colour_data = 24'b010100110011100001000111;
		12'b000001000000: colour_data = 24'b010100110011100001000111;
		12'b000001000001: colour_data = 24'b010100110011100001000111;
		12'b000001000010: colour_data = 24'b010100110011100001000111;
		12'b000001000011: colour_data = 24'b010100110011100001000111;
		12'b000001000100: colour_data = 24'b010100110011100001000111;
		12'b000001000101: colour_data = 24'b010100110011100001000111;
		12'b000001000110: colour_data = 24'b010100110011100001000111;
		12'b000001000111: colour_data = 24'b010100110011100001000111;
		12'b000001001000: colour_data = 24'b010100110011100001000111;
		12'b000001001001: colour_data = 24'b010100110011100001000111;
		12'b000001001010: colour_data = 24'b010100110011100001000111;
		12'b000001001011: colour_data = 24'b010100110011100001000111;
		12'b000001001100: colour_data = 24'b010100110011100001000111;
		12'b000001001101: colour_data = 24'b010100110011100001000111;
		12'b000001001110: colour_data = 24'b010100110011100001000111;
		12'b000001001111: colour_data = 24'b010100110011100001000111;
		12'b000001010000: colour_data = 24'b010100110011100001000111;
		12'b000001010001: colour_data = 24'b010100110011100001000111;
		12'b000001010010: colour_data = 24'b010100110011100001000111;
		12'b000001010011: colour_data = 24'b010100110011100001000111;
		12'b000001010100: colour_data = 24'b010100110011100001000111;
		12'b000001010101: colour_data = 24'b010100110011100001000111;
		12'b000001010110: colour_data = 24'b010100110011100001000111;
		12'b000001010111: colour_data = 24'b010100110011100001000111;
		12'b000001011000: colour_data = 24'b010100110011100001000111;
		12'b000001011001: colour_data = 24'b010100110011100001000111;
		12'b000001011010: colour_data = 24'b010100110011100001000111;
		12'b000001011011: colour_data = 24'b010100110011100001000111;
		12'b000001011100: colour_data = 24'b010100110011100001000111;
		12'b000001011101: colour_data = 24'b010100110011100001000111;
		12'b000001011110: colour_data = 24'b010100110011100001000111;
		12'b000001011111: colour_data = 24'b010100110011100001000111;
		12'b000001100000: colour_data = 24'b010100110011100001000111;
		12'b000001100001: colour_data = 24'b010100110011100001000111;
		12'b000001100010: colour_data = 24'b010100110011100001000111;
		12'b000001100011: colour_data = 24'b010100110011100001000111;
		12'b000001100100: colour_data = 24'b010100110011100001000111;
		12'b000001100101: colour_data = 24'b010100110011100001000111;
		12'b000001100110: colour_data = 24'b010100110011100001000111;
		12'b000001100111: colour_data = 24'b010100110011100001000111;
		12'b000001101000: colour_data = 24'b010100110011100001000111;
		12'b000001101001: colour_data = 24'b010100110011100001000111;
		12'b000001101010: colour_data = 24'b010100110011100001000111;
		12'b000001101011: colour_data = 24'b010100110011100001000111;
		12'b000001101100: colour_data = 24'b010100110011100001000111;
		12'b000001101101: colour_data = 24'b010100110011100001000111;
		12'b000001101110: colour_data = 24'b010100110011100001000111;
		12'b000001101111: colour_data = 24'b010100110011100001000111;
		12'b000001110000: colour_data = 24'b010100110011100001000111;
		12'b000001110001: colour_data = 24'b010100110011100001000111;
		12'b000001110010: colour_data = 24'b010100110011100001000111;
		12'b000001110011: colour_data = 24'b010100110011100001000111;
		12'b000001110100: colour_data = 24'b010100110011100001000111;
		12'b000001110101: colour_data = 24'b010100110011100001000111;
		12'b000001110110: colour_data = 24'b010100110011100001000111;
		12'b000001110111: colour_data = 24'b010100110011100001000111;
		12'b000001111000: colour_data = 24'b010100110011100001000111;
		12'b000001111001: colour_data = 24'b010100110011100001000111;
		12'b000001111010: colour_data = 24'b010100110011100001000111;
		12'b000001111011: colour_data = 24'b010100110011100001000111;
		12'b000001111100: colour_data = 24'b010100110011100001000111;
		12'b000001111101: colour_data = 24'b010100110011100001000111;
		12'b000001111110: colour_data = 24'b010100110011100001000111;
		12'b000001111111: colour_data = 24'b010100110011100001000111;
		12'b000010000000: colour_data = 24'b010100110011100001000111;
		12'b000010000001: colour_data = 24'b010100110011100001000111;
		12'b000010000010: colour_data = 24'b010100110011100001000111;
		12'b000010000011: colour_data = 24'b010100110011100001000111;
		12'b000010000100: colour_data = 24'b010100110011100001000111;
		12'b000010000101: colour_data = 24'b010100110011100001000111;
		12'b000010000110: colour_data = 24'b010100110011100001000111;
		12'b000010000111: colour_data = 24'b010100110011100001000111;
		12'b000010001000: colour_data = 24'b010100110011100001000111;
		12'b000010001001: colour_data = 24'b010100110011100001000111;
		12'b000010001010: colour_data = 24'b010100110011100001000111;
		12'b000010001011: colour_data = 24'b010100110011100001000111;

		12'b000100000000: colour_data = 24'b111001001111110010001011;
		12'b000100000001: colour_data = 24'b111001001111110010001011;
		12'b000100000010: colour_data = 24'b111001001111110010001011;
		12'b000100000011: colour_data = 24'b111001001111110010001011;
		12'b000100000100: colour_data = 24'b111001001111110010001011;
		12'b000100000101: colour_data = 24'b111001001111110010001011;
		12'b000100000110: colour_data = 24'b111001001111110010001011;
		12'b000100000111: colour_data = 24'b111001001111110010001011;
		12'b000100001000: colour_data = 24'b111001001111110010001011;
		12'b000100001001: colour_data = 24'b111001001111110010001011;
		12'b000100001010: colour_data = 24'b111001001111110010001011;
		12'b000100001011: colour_data = 24'b111001001111110010001011;
		12'b000100001100: colour_data = 24'b111001001111110010001011;
		12'b000100001101: colour_data = 24'b111001001111110010001011;
		12'b000100001110: colour_data = 24'b111001001111110010001011;
		12'b000100001111: colour_data = 24'b111001001111110010001011;
		12'b000100010000: colour_data = 24'b111001001111110010001011;
		12'b000100010001: colour_data = 24'b111001001111110010001011;
		12'b000100010010: colour_data = 24'b111001001111110010001011;
		12'b000100010011: colour_data = 24'b111001001111110010001011;
		12'b000100010100: colour_data = 24'b111001001111110010001011;
		12'b000100010101: colour_data = 24'b111001001111110010001011;
		12'b000100010110: colour_data = 24'b111001001111110010001011;
		12'b000100010111: colour_data = 24'b111001001111110010001011;
		12'b000100011000: colour_data = 24'b111001001111110010001011;
		12'b000100011001: colour_data = 24'b111001001111110010001011;
		12'b000100011010: colour_data = 24'b111001001111110010001011;
		12'b000100011011: colour_data = 24'b111001001111110010001011;
		12'b000100011100: colour_data = 24'b111001001111110010001011;
		12'b000100011101: colour_data = 24'b111001001111110010001011;
		12'b000100011110: colour_data = 24'b111001001111110010001011;
		12'b000100011111: colour_data = 24'b111001001111110010001011;
		12'b000100100000: colour_data = 24'b111001001111110010001011;
		12'b000100100001: colour_data = 24'b111001001111110010001011;
		12'b000100100010: colour_data = 24'b111001001111110010001011;
		12'b000100100011: colour_data = 24'b111001001111110010001011;
		12'b000100100100: colour_data = 24'b111001001111110010001011;
		12'b000100100101: colour_data = 24'b111001001111110010001011;
		12'b000100100110: colour_data = 24'b111001001111110010001011;
		12'b000100100111: colour_data = 24'b111001001111110010001011;
		12'b000100101000: colour_data = 24'b111001001111110010001011;
		12'b000100101001: colour_data = 24'b111001001111110010001011;
		12'b000100101010: colour_data = 24'b111001001111110010001011;
		12'b000100101011: colour_data = 24'b111001001111110010001011;
		12'b000100101100: colour_data = 24'b111001001111110010001011;
		12'b000100101101: colour_data = 24'b111001001111110010001011;
		12'b000100101110: colour_data = 24'b111001001111110010001011;
		12'b000100101111: colour_data = 24'b111001001111110010001011;
		12'b000100110000: colour_data = 24'b111001001111110010001011;
		12'b000100110001: colour_data = 24'b111001001111110010001011;
		12'b000100110010: colour_data = 24'b111001001111110010001011;
		12'b000100110011: colour_data = 24'b111001001111110010001011;
		12'b000100110100: colour_data = 24'b111001001111110010001011;
		12'b000100110101: colour_data = 24'b111001001111110010001011;
		12'b000100110110: colour_data = 24'b111001001111110010001011;
		12'b000100110111: colour_data = 24'b111001001111110010001011;
		12'b000100111000: colour_data = 24'b111001001111110010001011;
		12'b000100111001: colour_data = 24'b111001001111110010001011;
		12'b000100111010: colour_data = 24'b111001001111110010001011;
		12'b000100111011: colour_data = 24'b111001001111110010001011;
		12'b000100111100: colour_data = 24'b111001001111110010001011;
		12'b000100111101: colour_data = 24'b111001001111110010001011;
		12'b000100111110: colour_data = 24'b111001001111110010001011;
		12'b000100111111: colour_data = 24'b111001001111110010001011;
		12'b000101000000: colour_data = 24'b111001001111110010001011;
		12'b000101000001: colour_data = 24'b111001001111110010001011;
		12'b000101000010: colour_data = 24'b111001001111110010001011;
		12'b000101000011: colour_data = 24'b111001001111110010001011;
		12'b000101000100: colour_data = 24'b111001001111110010001011;
		12'b000101000101: colour_data = 24'b111001001111110010001011;
		12'b000101000110: colour_data = 24'b111001001111110010001011;
		12'b000101000111: colour_data = 24'b111001001111110010001011;
		12'b000101001000: colour_data = 24'b111001001111110010001011;
		12'b000101001001: colour_data = 24'b111001001111110010001011;
		12'b000101001010: colour_data = 24'b111001001111110010001011;
		12'b000101001011: colour_data = 24'b111001001111110010001011;
		12'b000101001100: colour_data = 24'b111001001111110010001011;
		12'b000101001101: colour_data = 24'b111001001111110010001011;
		12'b000101001110: colour_data = 24'b111001001111110010001011;
		12'b000101001111: colour_data = 24'b111001001111110010001011;
		12'b000101010000: colour_data = 24'b111001001111110010001011;
		12'b000101010001: colour_data = 24'b111001001111110010001011;
		12'b000101010010: colour_data = 24'b111001001111110010001011;
		12'b000101010011: colour_data = 24'b111001001111110010001011;
		12'b000101010100: colour_data = 24'b111001001111110010001011;
		12'b000101010101: colour_data = 24'b111001001111110010001011;
		12'b000101010110: colour_data = 24'b111001001111110010001011;
		12'b000101010111: colour_data = 24'b111001001111110010001011;
		12'b000101011000: colour_data = 24'b111001001111110010001011;
		12'b000101011001: colour_data = 24'b111001001111110010001011;
		12'b000101011010: colour_data = 24'b111001001111110010001011;
		12'b000101011011: colour_data = 24'b111001001111110010001011;
		12'b000101011100: colour_data = 24'b111001001111110010001011;
		12'b000101011101: colour_data = 24'b111001001111110010001011;
		12'b000101011110: colour_data = 24'b111001001111110010001011;
		12'b000101011111: colour_data = 24'b111001001111110010001011;
		12'b000101100000: colour_data = 24'b111001001111110010001011;
		12'b000101100001: colour_data = 24'b111001001111110010001011;
		12'b000101100010: colour_data = 24'b111001001111110010001011;
		12'b000101100011: colour_data = 24'b111001001111110010001011;
		12'b000101100100: colour_data = 24'b111001001111110010001011;
		12'b000101100101: colour_data = 24'b111001001111110010001011;
		12'b000101100110: colour_data = 24'b111001001111110010001011;
		12'b000101100111: colour_data = 24'b111001001111110010001011;
		12'b000101101000: colour_data = 24'b111001001111110010001011;
		12'b000101101001: colour_data = 24'b111001001111110010001011;
		12'b000101101010: colour_data = 24'b111001001111110010001011;
		12'b000101101011: colour_data = 24'b111001001111110010001011;
		12'b000101101100: colour_data = 24'b111001001111110010001011;
		12'b000101101101: colour_data = 24'b111001001111110010001011;
		12'b000101101110: colour_data = 24'b111001001111110010001011;
		12'b000101101111: colour_data = 24'b111001001111110010001011;
		12'b000101110000: colour_data = 24'b111001001111110010001011;
		12'b000101110001: colour_data = 24'b111001001111110010001011;
		12'b000101110010: colour_data = 24'b111001001111110010001011;
		12'b000101110011: colour_data = 24'b111001001111110010001011;
		12'b000101110100: colour_data = 24'b111001001111110010001011;
		12'b000101110101: colour_data = 24'b111001001111110010001011;
		12'b000101110110: colour_data = 24'b111001001111110010001011;
		12'b000101110111: colour_data = 24'b111001001111110010001011;
		12'b000101111000: colour_data = 24'b111001001111110010001011;
		12'b000101111001: colour_data = 24'b111001001111110010001011;
		12'b000101111010: colour_data = 24'b111001001111110010001011;
		12'b000101111011: colour_data = 24'b111001001111110010001011;
		12'b000101111100: colour_data = 24'b111001001111110010001011;
		12'b000101111101: colour_data = 24'b111001001111110010001011;
		12'b000101111110: colour_data = 24'b111001001111110010001011;
		12'b000101111111: colour_data = 24'b111001001111110010001011;
		12'b000110000000: colour_data = 24'b111001001111110010001011;
		12'b000110000001: colour_data = 24'b111001001111110010001011;
		12'b000110000010: colour_data = 24'b111001001111110010001011;
		12'b000110000011: colour_data = 24'b111001001111110010001011;
		12'b000110000100: colour_data = 24'b111001001111110010001011;
		12'b000110000101: colour_data = 24'b111001001111110010001011;
		12'b000110000110: colour_data = 24'b111001001111110010001011;
		12'b000110000111: colour_data = 24'b111001001111110010001011;
		12'b000110001000: colour_data = 24'b111001001111110010001011;
		12'b000110001001: colour_data = 24'b111001001111110010001011;
		12'b000110001010: colour_data = 24'b111001001111110010001011;
		12'b000110001011: colour_data = 24'b111001001111110010001011;

		12'b001000000000: colour_data = 24'b100111001110011001011001;
		12'b001000000001: colour_data = 24'b100111001110011001011001;
		12'b001000000010: colour_data = 24'b011100111011111100101110;
		12'b001000000011: colour_data = 24'b011100111011111100101110;
		12'b001000000100: colour_data = 24'b011100111011111100101110;
		12'b001000000101: colour_data = 24'b011100111011111100101110;
		12'b001000000110: colour_data = 24'b100111001110011001011001;
		12'b001000000111: colour_data = 24'b100111001110011001011001;
		12'b001000001000: colour_data = 24'b100111001110011001011001;
		12'b001000001001: colour_data = 24'b011100111011111100101110;
		12'b001000001010: colour_data = 24'b011100111011111100101110;
		12'b001000001011: colour_data = 24'b011100111011111100101110;
		12'b001000001100: colour_data = 24'b011100111011111100101110;
		12'b001000001101: colour_data = 24'b100111001110011001011001;
		12'b001000001110: colour_data = 24'b100111001110011001011001;
		12'b001000001111: colour_data = 24'b100111001110011001011001;
		12'b001000010000: colour_data = 24'b011100111011111100101110;
		12'b001000010001: colour_data = 24'b011100111011111100101110;
		12'b001000010010: colour_data = 24'b011100111011111100101110;
		12'b001000010011: colour_data = 24'b011100111011111100101110;
		12'b001000010100: colour_data = 24'b100111001110011001011001;
		12'b001000010101: colour_data = 24'b100111001110011001011001;
		12'b001000010110: colour_data = 24'b100111001110011001011001;
		12'b001000010111: colour_data = 24'b011100111011111100101110;
		12'b001000011000: colour_data = 24'b011100111011111100101110;
		12'b001000011001: colour_data = 24'b011100111011111100101110;
		12'b001000011010: colour_data = 24'b011100111011111100101110;
		12'b001000011011: colour_data = 24'b100111001110011001011001;
		12'b001000011100: colour_data = 24'b100111001110011001011001;
		12'b001000011101: colour_data = 24'b100111001110011001011001;
		12'b001000011110: colour_data = 24'b011100111011111100101110;
		12'b001000011111: colour_data = 24'b011100111011111100101110;
		12'b001000100000: colour_data = 24'b011100111011111100101110;
		12'b001000100001: colour_data = 24'b011100111011111100101110;
		12'b001000100010: colour_data = 24'b100111001110011001011001;
		12'b001000100011: colour_data = 24'b100111001110011001011001;
		12'b001000100100: colour_data = 24'b100111001110011001011001;
		12'b001000100101: colour_data = 24'b011100111011111100101110;
		12'b001000100110: colour_data = 24'b011100111011111100101110;
		12'b001000100111: colour_data = 24'b011100111011111100101110;
		12'b001000101000: colour_data = 24'b011100111011111100101110;
		12'b001000101001: colour_data = 24'b100111001110011001011001;
		12'b001000101010: colour_data = 24'b100111001110011001011001;
		12'b001000101011: colour_data = 24'b100111001110011001011001;
		12'b001000101100: colour_data = 24'b011100111011111100101110;
		12'b001000101101: colour_data = 24'b011100111011111100101110;
		12'b001000101110: colour_data = 24'b011100111011111100101110;
		12'b001000101111: colour_data = 24'b011100111011111100101110;
		12'b001000110000: colour_data = 24'b100111001110011001011001;
		12'b001000110001: colour_data = 24'b100111001110011001011001;
		12'b001000110010: colour_data = 24'b100111001110011001011001;
		12'b001000110011: colour_data = 24'b011100111011111100101110;
		12'b001000110100: colour_data = 24'b011100111011111100101110;
		12'b001000110101: colour_data = 24'b011100111011111100101110;
		12'b001000110110: colour_data = 24'b011100111011111100101110;
		12'b001000110111: colour_data = 24'b100111001110011001011001;
		12'b001000111000: colour_data = 24'b100111001110011001011001;
		12'b001000111001: colour_data = 24'b100111001110011001011001;
		12'b001000111010: colour_data = 24'b011100111011111100101110;
		12'b001000111011: colour_data = 24'b011100111011111100101110;
		12'b001000111100: colour_data = 24'b011100111011111100101110;
		12'b001000111101: colour_data = 24'b011100111011111100101110;
		12'b001000111110: colour_data = 24'b100111001110011001011001;
		12'b001000111111: colour_data = 24'b100111001110011001011001;
		12'b001001000000: colour_data = 24'b100111001110011001011001;
		12'b001001000001: colour_data = 24'b011100111011111100101110;
		12'b001001000010: colour_data = 24'b011100111011111100101110;
		12'b001001000011: colour_data = 24'b011100111011111100101110;
		12'b001001000100: colour_data = 24'b011100111011111100101110;
		12'b001001000101: colour_data = 24'b100111001110011001011001;
		12'b001001000110: colour_data = 24'b100111001110011001011001;
		12'b001001000111: colour_data = 24'b100111001110011001011001;
		12'b001001001000: colour_data = 24'b011100111011111100101110;
		12'b001001001001: colour_data = 24'b011100111011111100101110;
		12'b001001001010: colour_data = 24'b011100111011111100101110;
		12'b001001001011: colour_data = 24'b011100111011111100101110;
		12'b001001001100: colour_data = 24'b100111001110011001011001;
		12'b001001001101: colour_data = 24'b100111001110011001011001;
		12'b001001001110: colour_data = 24'b100111001110011001011001;
		12'b001001001111: colour_data = 24'b011100111011111100101110;
		12'b001001010000: colour_data = 24'b011100111011111100101110;
		12'b001001010001: colour_data = 24'b011100111011111100101110;
		12'b001001010010: colour_data = 24'b011100111011111100101110;
		12'b001001010011: colour_data = 24'b100111001110011001011001;
		12'b001001010100: colour_data = 24'b100111001110011001011001;
		12'b001001010101: colour_data = 24'b100111001110011001011001;
		12'b001001010110: colour_data = 24'b011100111011111100101110;
		12'b001001010111: colour_data = 24'b011100111011111100101110;
		12'b001001011000: colour_data = 24'b011100111011111100101110;
		12'b001001011001: colour_data = 24'b011100111011111100101110;
		12'b001001011010: colour_data = 24'b100111001110011001011001;
		12'b001001011011: colour_data = 24'b100111001110011001011001;
		12'b001001011100: colour_data = 24'b100111001110011001011001;
		12'b001001011101: colour_data = 24'b011100111011111100101110;
		12'b001001011110: colour_data = 24'b011100111011111100101110;
		12'b001001011111: colour_data = 24'b011100111011111100101110;
		12'b001001100000: colour_data = 24'b011100111011111100101110;
		12'b001001100001: colour_data = 24'b100111001110011001011001;
		12'b001001100010: colour_data = 24'b100111001110011001011001;
		12'b001001100011: colour_data = 24'b100111001110011001011001;
		12'b001001100100: colour_data = 24'b011100111011111100101110;
		12'b001001100101: colour_data = 24'b011100111011111100101110;
		12'b001001100110: colour_data = 24'b011100111011111100101110;
		12'b001001100111: colour_data = 24'b011100111011111100101110;
		12'b001001101000: colour_data = 24'b100111001110011001011001;
		12'b001001101001: colour_data = 24'b100111001110011001011001;
		12'b001001101010: colour_data = 24'b100111001110011001011001;
		12'b001001101011: colour_data = 24'b011100111011111100101110;
		12'b001001101100: colour_data = 24'b011100111011111100101110;
		12'b001001101101: colour_data = 24'b011100111011111100101110;
		12'b001001101110: colour_data = 24'b011100111011111100101110;
		12'b001001101111: colour_data = 24'b100111001110011001011001;
		12'b001001110000: colour_data = 24'b100111001110011001011001;
		12'b001001110001: colour_data = 24'b100111001110011001011001;
		12'b001001110010: colour_data = 24'b011100111011111100101110;
		12'b001001110011: colour_data = 24'b011100111011111100101110;
		12'b001001110100: colour_data = 24'b011100111011111100101110;
		12'b001001110101: colour_data = 24'b011100111011111100101110;
		12'b001001110110: colour_data = 24'b100111001110011001011001;
		12'b001001110111: colour_data = 24'b100111001110011001011001;
		12'b001001111000: colour_data = 24'b100111001110011001011001;
		12'b001001111001: colour_data = 24'b011100111011111100101110;
		12'b001001111010: colour_data = 24'b011100111011111100101110;
		12'b001001111011: colour_data = 24'b011100111011111100101110;
		12'b001001111100: colour_data = 24'b011100111011111100101110;
		12'b001001111101: colour_data = 24'b100111001110011001011001;
		12'b001001111110: colour_data = 24'b100111001110011001011001;
		12'b001001111111: colour_data = 24'b100111001110011001011001;
		12'b001010000000: colour_data = 24'b011100111011111100101110;
		12'b001010000001: colour_data = 24'b011100111011111100101110;
		12'b001010000010: colour_data = 24'b011100111011111100101110;
		12'b001010000011: colour_data = 24'b011100111011111100101110;
		12'b001010000100: colour_data = 24'b100111001110011001011001;
		12'b001010000101: colour_data = 24'b100111001110011001011001;
		12'b001010000110: colour_data = 24'b100111001110011001011001;
		12'b001010000111: colour_data = 24'b011100111011111100101110;
		12'b001010001000: colour_data = 24'b011100111011111100101110;
		12'b001010001001: colour_data = 24'b011100111011111100101110;
		12'b001010001010: colour_data = 24'b011100111011111100101110;
		12'b001010001011: colour_data = 24'b100111001110011001011001;

		12'b001100000000: colour_data = 24'b100111001110011001011001;
		12'b001100000001: colour_data = 24'b011100111011111100101110;
		12'b001100000010: colour_data = 24'b011100111011111100101110;
		12'b001100000011: colour_data = 24'b011100111011111100101110;
		12'b001100000100: colour_data = 24'b011100111011111100101110;
		12'b001100000101: colour_data = 24'b100111001110011001011001;
		12'b001100000110: colour_data = 24'b100111001110011001011001;
		12'b001100000111: colour_data = 24'b100111001110011001011001;
		12'b001100001000: colour_data = 24'b011100111011111100101110;
		12'b001100001001: colour_data = 24'b011100111011111100101110;
		12'b001100001010: colour_data = 24'b011100111011111100101110;
		12'b001100001011: colour_data = 24'b011100111011111100101110;
		12'b001100001100: colour_data = 24'b100111001110011001011001;
		12'b001100001101: colour_data = 24'b100111001110011001011001;
		12'b001100001110: colour_data = 24'b100111001110011001011001;
		12'b001100001111: colour_data = 24'b011100111011111100101110;
		12'b001100010000: colour_data = 24'b011100111011111100101110;
		12'b001100010001: colour_data = 24'b011100111011111100101110;
		12'b001100010010: colour_data = 24'b011100111011111100101110;
		12'b001100010011: colour_data = 24'b100111001110011001011001;
		12'b001100010100: colour_data = 24'b100111001110011001011001;
		12'b001100010101: colour_data = 24'b100111001110011001011001;
		12'b001100010110: colour_data = 24'b011100111011111100101110;
		12'b001100010111: colour_data = 24'b011100111011111100101110;
		12'b001100011000: colour_data = 24'b011100111011111100101110;
		12'b001100011001: colour_data = 24'b011100111011111100101110;
		12'b001100011010: colour_data = 24'b100111001110011001011001;
		12'b001100011011: colour_data = 24'b100111001110011001011001;
		12'b001100011100: colour_data = 24'b100111001110011001011001;
		12'b001100011101: colour_data = 24'b011100111011111100101110;
		12'b001100011110: colour_data = 24'b011100111011111100101110;
		12'b001100011111: colour_data = 24'b011100111011111100101110;
		12'b001100100000: colour_data = 24'b011100111011111100101110;
		12'b001100100001: colour_data = 24'b100111001110011001011001;
		12'b001100100010: colour_data = 24'b100111001110011001011001;
		12'b001100100011: colour_data = 24'b100111001110011001011001;
		12'b001100100100: colour_data = 24'b011100111011111100101110;
		12'b001100100101: colour_data = 24'b011100111011111100101110;
		12'b001100100110: colour_data = 24'b011100111011111100101110;
		12'b001100100111: colour_data = 24'b011100111011111100101110;
		12'b001100101000: colour_data = 24'b100111001110011001011001;
		12'b001100101001: colour_data = 24'b100111001110011001011001;
		12'b001100101010: colour_data = 24'b100111001110011001011001;
		12'b001100101011: colour_data = 24'b011100111011111100101110;
		12'b001100101100: colour_data = 24'b011100111011111100101110;
		12'b001100101101: colour_data = 24'b011100111011111100101110;
		12'b001100101110: colour_data = 24'b011100111011111100101110;
		12'b001100101111: colour_data = 24'b100111001110011001011001;
		12'b001100110000: colour_data = 24'b100111001110011001011001;
		12'b001100110001: colour_data = 24'b100111001110011001011001;
		12'b001100110010: colour_data = 24'b011100111011111100101110;
		12'b001100110011: colour_data = 24'b011100111011111100101110;
		12'b001100110100: colour_data = 24'b011100111011111100101110;
		12'b001100110101: colour_data = 24'b011100111011111100101110;
		12'b001100110110: colour_data = 24'b100111001110011001011001;
		12'b001100110111: colour_data = 24'b100111001110011001011001;
		12'b001100111000: colour_data = 24'b100111001110011001011001;
		12'b001100111001: colour_data = 24'b011100111011111100101110;
		12'b001100111010: colour_data = 24'b011100111011111100101110;
		12'b001100111011: colour_data = 24'b011100111011111100101110;
		12'b001100111100: colour_data = 24'b011100111011111100101110;
		12'b001100111101: colour_data = 24'b100111001110011001011001;
		12'b001100111110: colour_data = 24'b100111001110011001011001;
		12'b001100111111: colour_data = 24'b100111001110011001011001;
		12'b001101000000: colour_data = 24'b011100111011111100101110;
		12'b001101000001: colour_data = 24'b011100111011111100101110;
		12'b001101000010: colour_data = 24'b011100111011111100101110;
		12'b001101000011: colour_data = 24'b011100111011111100101110;
		12'b001101000100: colour_data = 24'b100111001110011001011001;
		12'b001101000101: colour_data = 24'b100111001110011001011001;
		12'b001101000110: colour_data = 24'b100111001110011001011001;
		12'b001101000111: colour_data = 24'b011100111011111100101110;
		12'b001101001000: colour_data = 24'b011100111011111100101110;
		12'b001101001001: colour_data = 24'b011100111011111100101110;
		12'b001101001010: colour_data = 24'b011100111011111100101110;
		12'b001101001011: colour_data = 24'b100111001110011001011001;
		12'b001101001100: colour_data = 24'b100111001110011001011001;
		12'b001101001101: colour_data = 24'b100111001110011001011001;
		12'b001101001110: colour_data = 24'b011100111011111100101110;
		12'b001101001111: colour_data = 24'b011100111011111100101110;
		12'b001101010000: colour_data = 24'b011100111011111100101110;
		12'b001101010001: colour_data = 24'b011100111011111100101110;
		12'b001101010010: colour_data = 24'b100111001110011001011001;
		12'b001101010011: colour_data = 24'b100111001110011001011001;
		12'b001101010100: colour_data = 24'b100111001110011001011001;
		12'b001101010101: colour_data = 24'b011100111011111100101110;
		12'b001101010110: colour_data = 24'b011100111011111100101110;
		12'b001101010111: colour_data = 24'b011100111011111100101110;
		12'b001101011000: colour_data = 24'b011100111011111100101110;
		12'b001101011001: colour_data = 24'b100111001110011001011001;
		12'b001101011010: colour_data = 24'b100111001110011001011001;
		12'b001101011011: colour_data = 24'b100111001110011001011001;
		12'b001101011100: colour_data = 24'b011100111011111100101110;
		12'b001101011101: colour_data = 24'b011100111011111100101110;
		12'b001101011110: colour_data = 24'b011100111011111100101110;
		12'b001101011111: colour_data = 24'b011100111011111100101110;
		12'b001101100000: colour_data = 24'b100111001110011001011001;
		12'b001101100001: colour_data = 24'b100111001110011001011001;
		12'b001101100010: colour_data = 24'b100111001110011001011001;
		12'b001101100011: colour_data = 24'b011100111011111100101110;
		12'b001101100100: colour_data = 24'b011100111011111100101110;
		12'b001101100101: colour_data = 24'b011100111011111100101110;
		12'b001101100110: colour_data = 24'b011100111011111100101110;
		12'b001101100111: colour_data = 24'b100111001110011001011001;
		12'b001101101000: colour_data = 24'b100111001110011001011001;
		12'b001101101001: colour_data = 24'b100111001110011001011001;
		12'b001101101010: colour_data = 24'b011100111011111100101110;
		12'b001101101011: colour_data = 24'b011100111011111100101110;
		12'b001101101100: colour_data = 24'b011100111011111100101110;
		12'b001101101101: colour_data = 24'b011100111011111100101110;
		12'b001101101110: colour_data = 24'b100111001110011001011001;
		12'b001101101111: colour_data = 24'b100111001110011001011001;
		12'b001101110000: colour_data = 24'b100111001110011001011001;
		12'b001101110001: colour_data = 24'b011100111011111100101110;
		12'b001101110010: colour_data = 24'b011100111011111100101110;
		12'b001101110011: colour_data = 24'b011100111011111100101110;
		12'b001101110100: colour_data = 24'b011100111011111100101110;
		12'b001101110101: colour_data = 24'b100111001110011001011001;
		12'b001101110110: colour_data = 24'b100111001110011001011001;
		12'b001101110111: colour_data = 24'b100111001110011001011001;
		12'b001101111000: colour_data = 24'b011100111011111100101110;
		12'b001101111001: colour_data = 24'b011100111011111100101110;
		12'b001101111010: colour_data = 24'b011100111011111100101110;
		12'b001101111011: colour_data = 24'b011100111011111100101110;
		12'b001101111100: colour_data = 24'b100111001110011001011001;
		12'b001101111101: colour_data = 24'b100111001110011001011001;
		12'b001101111110: colour_data = 24'b100111001110011001011001;
		12'b001101111111: colour_data = 24'b011100111011111100101110;
		12'b001110000000: colour_data = 24'b011100111011111100101110;
		12'b001110000001: colour_data = 24'b011100111011111100101110;
		12'b001110000010: colour_data = 24'b011100111011111100101110;
		12'b001110000011: colour_data = 24'b100111001110011001011001;
		12'b001110000100: colour_data = 24'b100111001110011001011001;
		12'b001110000101: colour_data = 24'b100111001110011001011001;
		12'b001110000110: colour_data = 24'b011100111011111100101110;
		12'b001110000111: colour_data = 24'b011100111011111100101110;
		12'b001110001000: colour_data = 24'b011100111011111100101110;
		12'b001110001001: colour_data = 24'b011100111011111100101110;
		12'b001110001010: colour_data = 24'b100111001110011001011001;
		12'b001110001011: colour_data = 24'b100111001110011001011001;

		12'b010000000000: colour_data = 24'b011100111011111100101110;
		12'b010000000001: colour_data = 24'b011100111011111100101110;
		12'b010000000010: colour_data = 24'b011100111011111100101110;
		12'b010000000011: colour_data = 24'b011100111011111100101110;
		12'b010000000100: colour_data = 24'b100111001110011001011001;
		12'b010000000101: colour_data = 24'b100111001110011001011001;
		12'b010000000110: colour_data = 24'b100111001110011001011001;
		12'b010000000111: colour_data = 24'b011100111011111100101110;
		12'b010000001000: colour_data = 24'b011100111011111100101110;
		12'b010000001001: colour_data = 24'b011100111011111100101110;
		12'b010000001010: colour_data = 24'b011100111011111100101110;
		12'b010000001011: colour_data = 24'b100111001110011001011001;
		12'b010000001100: colour_data = 24'b100111001110011001011001;
		12'b010000001101: colour_data = 24'b100111001110011001011001;
		12'b010000001110: colour_data = 24'b011100111011111100101110;
		12'b010000001111: colour_data = 24'b011100111011111100101110;
		12'b010000010000: colour_data = 24'b011100111011111100101110;
		12'b010000010001: colour_data = 24'b011100111011111100101110;
		12'b010000010010: colour_data = 24'b100111001110011001011001;
		12'b010000010011: colour_data = 24'b100111001110011001011001;
		12'b010000010100: colour_data = 24'b100111001110011001011001;
		12'b010000010101: colour_data = 24'b011100111011111100101110;
		12'b010000010110: colour_data = 24'b011100111011111100101110;
		12'b010000010111: colour_data = 24'b011100111011111100101110;
		12'b010000011000: colour_data = 24'b011100111011111100101110;
		12'b010000011001: colour_data = 24'b100111001110011001011001;
		12'b010000011010: colour_data = 24'b100111001110011001011001;
		12'b010000011011: colour_data = 24'b100111001110011001011001;
		12'b010000011100: colour_data = 24'b011100111011111100101110;
		12'b010000011101: colour_data = 24'b011100111011111100101110;
		12'b010000011110: colour_data = 24'b011100111011111100101110;
		12'b010000011111: colour_data = 24'b011100111011111100101110;
		12'b010000100000: colour_data = 24'b100111001110011001011001;
		12'b010000100001: colour_data = 24'b100111001110011001011001;
		12'b010000100010: colour_data = 24'b100111001110011001011001;
		12'b010000100011: colour_data = 24'b011100111011111100101110;
		12'b010000100100: colour_data = 24'b011100111011111100101110;
		12'b010000100101: colour_data = 24'b011100111011111100101110;
		12'b010000100110: colour_data = 24'b011100111011111100101110;
		12'b010000100111: colour_data = 24'b100111001110011001011001;
		12'b010000101000: colour_data = 24'b100111001110011001011001;
		12'b010000101001: colour_data = 24'b100111001110011001011001;
		12'b010000101010: colour_data = 24'b011100111011111100101110;
		12'b010000101011: colour_data = 24'b011100111011111100101110;
		12'b010000101100: colour_data = 24'b011100111011111100101110;
		12'b010000101101: colour_data = 24'b011100111011111100101110;
		12'b010000101110: colour_data = 24'b100111001110011001011001;
		12'b010000101111: colour_data = 24'b100111001110011001011001;
		12'b010000110000: colour_data = 24'b100111001110011001011001;
		12'b010000110001: colour_data = 24'b011100111011111100101110;
		12'b010000110010: colour_data = 24'b011100111011111100101110;
		12'b010000110011: colour_data = 24'b011100111011111100101110;
		12'b010000110100: colour_data = 24'b011100111011111100101110;
		12'b010000110101: colour_data = 24'b100111001110011001011001;
		12'b010000110110: colour_data = 24'b100111001110011001011001;
		12'b010000110111: colour_data = 24'b100111001110011001011001;
		12'b010000111000: colour_data = 24'b011100111011111100101110;
		12'b010000111001: colour_data = 24'b011100111011111100101110;
		12'b010000111010: colour_data = 24'b011100111011111100101110;
		12'b010000111011: colour_data = 24'b011100111011111100101110;
		12'b010000111100: colour_data = 24'b100111001110011001011001;
		12'b010000111101: colour_data = 24'b100111001110011001011001;
		12'b010000111110: colour_data = 24'b100111001110011001011001;
		12'b010000111111: colour_data = 24'b011100111011111100101110;
		12'b010001000000: colour_data = 24'b011100111011111100101110;
		12'b010001000001: colour_data = 24'b011100111011111100101110;
		12'b010001000010: colour_data = 24'b011100111011111100101110;
		12'b010001000011: colour_data = 24'b100111001110011001011001;
		12'b010001000100: colour_data = 24'b100111001110011001011001;
		12'b010001000101: colour_data = 24'b100111001110011001011001;
		12'b010001000110: colour_data = 24'b011100111011111100101110;
		12'b010001000111: colour_data = 24'b011100111011111100101110;
		12'b010001001000: colour_data = 24'b011100111011111100101110;
		12'b010001001001: colour_data = 24'b011100111011111100101110;
		12'b010001001010: colour_data = 24'b100111001110011001011001;
		12'b010001001011: colour_data = 24'b100111001110011001011001;
		12'b010001001100: colour_data = 24'b100111001110011001011001;
		12'b010001001101: colour_data = 24'b011100111011111100101110;
		12'b010001001110: colour_data = 24'b011100111011111100101110;
		12'b010001001111: colour_data = 24'b011100111011111100101110;
		12'b010001010000: colour_data = 24'b011100111011111100101110;
		12'b010001010001: colour_data = 24'b100111001110011001011001;
		12'b010001010010: colour_data = 24'b100111001110011001011001;
		12'b010001010011: colour_data = 24'b100111001110011001011001;
		12'b010001010100: colour_data = 24'b011100111011111100101110;
		12'b010001010101: colour_data = 24'b011100111011111100101110;
		12'b010001010110: colour_data = 24'b011100111011111100101110;
		12'b010001010111: colour_data = 24'b011100111011111100101110;
		12'b010001011000: colour_data = 24'b100111001110011001011001;
		12'b010001011001: colour_data = 24'b100111001110011001011001;
		12'b010001011010: colour_data = 24'b100111001110011001011001;
		12'b010001011011: colour_data = 24'b011100111011111100101110;
		12'b010001011100: colour_data = 24'b011100111011111100101110;
		12'b010001011101: colour_data = 24'b011100111011111100101110;
		12'b010001011110: colour_data = 24'b011100111011111100101110;
		12'b010001011111: colour_data = 24'b100111001110011001011001;
		12'b010001100000: colour_data = 24'b100111001110011001011001;
		12'b010001100001: colour_data = 24'b100111001110011001011001;
		12'b010001100010: colour_data = 24'b011100111011111100101110;
		12'b010001100011: colour_data = 24'b011100111011111100101110;
		12'b010001100100: colour_data = 24'b011100111011111100101110;
		12'b010001100101: colour_data = 24'b011100111011111100101110;
		12'b010001100110: colour_data = 24'b100111001110011001011001;
		12'b010001100111: colour_data = 24'b100111001110011001011001;
		12'b010001101000: colour_data = 24'b100111001110011001011001;
		12'b010001101001: colour_data = 24'b011100111011111100101110;
		12'b010001101010: colour_data = 24'b011100111011111100101110;
		12'b010001101011: colour_data = 24'b011100111011111100101110;
		12'b010001101100: colour_data = 24'b011100111011111100101110;
		12'b010001101101: colour_data = 24'b100111001110011001011001;
		12'b010001101110: colour_data = 24'b100111001110011001011001;
		12'b010001101111: colour_data = 24'b100111001110011001011001;
		12'b010001110000: colour_data = 24'b011100111011111100101110;
		12'b010001110001: colour_data = 24'b011100111011111100101110;
		12'b010001110010: colour_data = 24'b011100111011111100101110;
		12'b010001110011: colour_data = 24'b011100111011111100101110;
		12'b010001110100: colour_data = 24'b100111001110011001011001;
		12'b010001110101: colour_data = 24'b100111001110011001011001;
		12'b010001110110: colour_data = 24'b100111001110011001011001;
		12'b010001110111: colour_data = 24'b011100111011111100101110;
		12'b010001111000: colour_data = 24'b011100111011111100101110;
		12'b010001111001: colour_data = 24'b011100111011111100101110;
		12'b010001111010: colour_data = 24'b011100111011111100101110;
		12'b010001111011: colour_data = 24'b100111001110011001011001;
		12'b010001111100: colour_data = 24'b100111001110011001011001;
		12'b010001111101: colour_data = 24'b100111001110011001011001;
		12'b010001111110: colour_data = 24'b011100111011111100101110;
		12'b010001111111: colour_data = 24'b011100111011111100101110;
		12'b010010000000: colour_data = 24'b011100111011111100101110;
		12'b010010000001: colour_data = 24'b011100111011111100101110;
		12'b010010000010: colour_data = 24'b100111001110011001011001;
		12'b010010000011: colour_data = 24'b100111001110011001011001;
		12'b010010000100: colour_data = 24'b100111001110011001011001;
		12'b010010000101: colour_data = 24'b011100111011111100101110;
		12'b010010000110: colour_data = 24'b011100111011111100101110;
		12'b010010000111: colour_data = 24'b011100111011111100101110;
		12'b010010001000: colour_data = 24'b011100111011111100101110;
		12'b010010001001: colour_data = 24'b100111001110011001011001;
		12'b010010001010: colour_data = 24'b100111001110011001011001;
		12'b010010001011: colour_data = 24'b100111001110011001011001;

		12'b010100000000: colour_data = 24'b010101011000000000100010;
		12'b010100000001: colour_data = 24'b010101011000000000100010;
		12'b010100000010: colour_data = 24'b010101011000000000100010;
		12'b010100000011: colour_data = 24'b010101011000000000100010;
		12'b010100000100: colour_data = 24'b010101011000000000100010;
		12'b010100000101: colour_data = 24'b010101011000000000100010;
		12'b010100000110: colour_data = 24'b010101011000000000100010;
		12'b010100000111: colour_data = 24'b010101011000000000100010;
		12'b010100001000: colour_data = 24'b010101011000000000100010;
		12'b010100001001: colour_data = 24'b010101011000000000100010;
		12'b010100001010: colour_data = 24'b010101011000000000100010;
		12'b010100001011: colour_data = 24'b010101011000000000100010;
		12'b010100001100: colour_data = 24'b010101011000000000100010;
		12'b010100001101: colour_data = 24'b010101011000000000100010;
		12'b010100001110: colour_data = 24'b010101011000000000100010;
		12'b010100001111: colour_data = 24'b010101011000000000100010;
		12'b010100010000: colour_data = 24'b010101011000000000100010;
		12'b010100010001: colour_data = 24'b010101011000000000100010;
		12'b010100010010: colour_data = 24'b010101011000000000100010;
		12'b010100010011: colour_data = 24'b010101011000000000100010;
		12'b010100010100: colour_data = 24'b010101011000000000100010;
		12'b010100010101: colour_data = 24'b010101011000000000100010;
		12'b010100010110: colour_data = 24'b010101011000000000100010;
		12'b010100010111: colour_data = 24'b010101011000000000100010;
		12'b010100011000: colour_data = 24'b010101011000000000100010;
		12'b010100011001: colour_data = 24'b010101011000000000100010;
		12'b010100011010: colour_data = 24'b010101011000000000100010;
		12'b010100011011: colour_data = 24'b010101011000000000100010;
		12'b010100011100: colour_data = 24'b010101011000000000100010;
		12'b010100011101: colour_data = 24'b010101011000000000100010;
		12'b010100011110: colour_data = 24'b010101011000000000100010;
		12'b010100011111: colour_data = 24'b010101011000000000100010;
		12'b010100100000: colour_data = 24'b010101011000000000100010;
		12'b010100100001: colour_data = 24'b010101011000000000100010;
		12'b010100100010: colour_data = 24'b010101011000000000100010;
		12'b010100100011: colour_data = 24'b010101011000000000100010;
		12'b010100100100: colour_data = 24'b010101011000000000100010;
		12'b010100100101: colour_data = 24'b010101011000000000100010;
		12'b010100100110: colour_data = 24'b010101011000000000100010;
		12'b010100100111: colour_data = 24'b010101011000000000100010;
		12'b010100101000: colour_data = 24'b010101011000000000100010;
		12'b010100101001: colour_data = 24'b010101011000000000100010;
		12'b010100101010: colour_data = 24'b010101011000000000100010;
		12'b010100101011: colour_data = 24'b010101011000000000100010;
		12'b010100101100: colour_data = 24'b010101011000000000100010;
		12'b010100101101: colour_data = 24'b010101011000000000100010;
		12'b010100101110: colour_data = 24'b010101011000000000100010;
		12'b010100101111: colour_data = 24'b010101011000000000100010;
		12'b010100110000: colour_data = 24'b010101011000000000100010;
		12'b010100110001: colour_data = 24'b010101011000000000100010;
		12'b010100110010: colour_data = 24'b010101011000000000100010;
		12'b010100110011: colour_data = 24'b010101011000000000100010;
		12'b010100110100: colour_data = 24'b010101011000000000100010;
		12'b010100110101: colour_data = 24'b010101011000000000100010;
		12'b010100110110: colour_data = 24'b010101011000000000100010;
		12'b010100110111: colour_data = 24'b010101011000000000100010;
		12'b010100111000: colour_data = 24'b010101011000000000100010;
		12'b010100111001: colour_data = 24'b010101011000000000100010;
		12'b010100111010: colour_data = 24'b010101011000000000100010;
		12'b010100111011: colour_data = 24'b010101011000000000100010;
		12'b010100111100: colour_data = 24'b010101011000000000100010;
		12'b010100111101: colour_data = 24'b010101011000000000100010;
		12'b010100111110: colour_data = 24'b010101011000000000100010;
		12'b010100111111: colour_data = 24'b010101011000000000100010;
		12'b010101000000: colour_data = 24'b010101011000000000100010;
		12'b010101000001: colour_data = 24'b010101011000000000100010;
		12'b010101000010: colour_data = 24'b010101011000000000100010;
		12'b010101000011: colour_data = 24'b010101011000000000100010;
		12'b010101000100: colour_data = 24'b010101011000000000100010;
		12'b010101000101: colour_data = 24'b010101011000000000100010;
		12'b010101000110: colour_data = 24'b010101011000000000100010;
		12'b010101000111: colour_data = 24'b010101011000000000100010;
		12'b010101001000: colour_data = 24'b010101011000000000100010;
		12'b010101001001: colour_data = 24'b010101011000000000100010;
		12'b010101001010: colour_data = 24'b010101011000000000100010;
		12'b010101001011: colour_data = 24'b010101011000000000100010;
		12'b010101001100: colour_data = 24'b010101011000000000100010;
		12'b010101001101: colour_data = 24'b010101011000000000100010;
		12'b010101001110: colour_data = 24'b010101011000000000100010;
		12'b010101001111: colour_data = 24'b010101011000000000100010;
		12'b010101010000: colour_data = 24'b010101011000000000100010;
		12'b010101010001: colour_data = 24'b010101011000000000100010;
		12'b010101010010: colour_data = 24'b010101011000000000100010;
		12'b010101010011: colour_data = 24'b010101011000000000100010;
		12'b010101010100: colour_data = 24'b010101011000000000100010;
		12'b010101010101: colour_data = 24'b010101011000000000100010;
		12'b010101010110: colour_data = 24'b010101011000000000100010;
		12'b010101010111: colour_data = 24'b010101011000000000100010;
		12'b010101011000: colour_data = 24'b010101011000000000100010;
		12'b010101011001: colour_data = 24'b010101011000000000100010;
		12'b010101011010: colour_data = 24'b010101011000000000100010;
		12'b010101011011: colour_data = 24'b010101011000000000100010;
		12'b010101011100: colour_data = 24'b010101011000000000100010;
		12'b010101011101: colour_data = 24'b010101011000000000100010;
		12'b010101011110: colour_data = 24'b010101011000000000100010;
		12'b010101011111: colour_data = 24'b010101011000000000100010;
		12'b010101100000: colour_data = 24'b010101011000000000100010;
		12'b010101100001: colour_data = 24'b010101011000000000100010;
		12'b010101100010: colour_data = 24'b010101011000000000100010;
		12'b010101100011: colour_data = 24'b010101011000000000100010;
		12'b010101100100: colour_data = 24'b010101011000000000100010;
		12'b010101100101: colour_data = 24'b010101011000000000100010;
		12'b010101100110: colour_data = 24'b010101011000000000100010;
		12'b010101100111: colour_data = 24'b010101011000000000100010;
		12'b010101101000: colour_data = 24'b010101011000000000100010;
		12'b010101101001: colour_data = 24'b010101011000000000100010;
		12'b010101101010: colour_data = 24'b010101011000000000100010;
		12'b010101101011: colour_data = 24'b010101011000000000100010;
		12'b010101101100: colour_data = 24'b010101011000000000100010;
		12'b010101101101: colour_data = 24'b010101011000000000100010;
		12'b010101101110: colour_data = 24'b010101011000000000100010;
		12'b010101101111: colour_data = 24'b010101011000000000100010;
		12'b010101110000: colour_data = 24'b010101011000000000100010;
		12'b010101110001: colour_data = 24'b010101011000000000100010;
		12'b010101110010: colour_data = 24'b010101011000000000100010;
		12'b010101110011: colour_data = 24'b010101011000000000100010;
		12'b010101110100: colour_data = 24'b010101011000000000100010;
		12'b010101110101: colour_data = 24'b010101011000000000100010;
		12'b010101110110: colour_data = 24'b010101011000000000100010;
		12'b010101110111: colour_data = 24'b010101011000000000100010;
		12'b010101111000: colour_data = 24'b010101011000000000100010;
		12'b010101111001: colour_data = 24'b010101011000000000100010;
		12'b010101111010: colour_data = 24'b010101011000000000100010;
		12'b010101111011: colour_data = 24'b010101011000000000100010;
		12'b010101111100: colour_data = 24'b010101011000000000100010;
		12'b010101111101: colour_data = 24'b010101011000000000100010;
		12'b010101111110: colour_data = 24'b010101011000000000100010;
		12'b010101111111: colour_data = 24'b010101011000000000100010;
		12'b010110000000: colour_data = 24'b010101011000000000100010;
		12'b010110000001: colour_data = 24'b010101011000000000100010;
		12'b010110000010: colour_data = 24'b010101011000000000100010;
		12'b010110000011: colour_data = 24'b010101011000000000100010;
		12'b010110000100: colour_data = 24'b010101011000000000100010;
		12'b010110000101: colour_data = 24'b010101011000000000100010;
		12'b010110000110: colour_data = 24'b010101011000000000100010;
		12'b010110000111: colour_data = 24'b010101011000000000100010;
		12'b010110001000: colour_data = 24'b010101011000000000100010;
		12'b010110001001: colour_data = 24'b010101011000000000100010;
		12'b010110001010: colour_data = 24'b010101011000000000100010;
		12'b010110001011: colour_data = 24'b010101011000000000100010;

		12'b011000000000: colour_data = 24'b110101111010100001001100;
		12'b011000000001: colour_data = 24'b110101111010100001001100;
		12'b011000000010: colour_data = 24'b110101111010100001001100;
		12'b011000000011: colour_data = 24'b110101111010100001001100;
		12'b011000000100: colour_data = 24'b110101111010100001001100;
		12'b011000000101: colour_data = 24'b110101111010100001001100;
		12'b011000000110: colour_data = 24'b110101111010100001001100;
		12'b011000000111: colour_data = 24'b110101111010100001001100;
		12'b011000001000: colour_data = 24'b110101111010100001001100;
		12'b011000001001: colour_data = 24'b110101111010100001001100;
		12'b011000001010: colour_data = 24'b110101111010100001001100;
		12'b011000001011: colour_data = 24'b110101111010100001001100;
		12'b011000001100: colour_data = 24'b110101111010100001001100;
		12'b011000001101: colour_data = 24'b110101111010100001001100;
		12'b011000001110: colour_data = 24'b110101111010100001001100;
		12'b011000001111: colour_data = 24'b110101111010100001001100;
		12'b011000010000: colour_data = 24'b110101111010100001001100;
		12'b011000010001: colour_data = 24'b110101111010100001001100;
		12'b011000010010: colour_data = 24'b110101111010100001001100;
		12'b011000010011: colour_data = 24'b110101111010100001001100;
		12'b011000010100: colour_data = 24'b110101111010100001001100;
		12'b011000010101: colour_data = 24'b110101111010100001001100;
		12'b011000010110: colour_data = 24'b110101111010100001001100;
		12'b011000010111: colour_data = 24'b110101111010100001001100;
		12'b011000011000: colour_data = 24'b110101111010100001001100;
		12'b011000011001: colour_data = 24'b110101111010100001001100;
		12'b011000011010: colour_data = 24'b110101111010100001001100;
		12'b011000011011: colour_data = 24'b110101111010100001001100;
		12'b011000011100: colour_data = 24'b110101111010100001001100;
		12'b011000011101: colour_data = 24'b110101111010100001001100;
		12'b011000011110: colour_data = 24'b110101111010100001001100;
		12'b011000011111: colour_data = 24'b110101111010100001001100;
		12'b011000100000: colour_data = 24'b110101111010100001001100;
		12'b011000100001: colour_data = 24'b110101111010100001001100;
		12'b011000100010: colour_data = 24'b110101111010100001001100;
		12'b011000100011: colour_data = 24'b110101111010100001001100;
		12'b011000100100: colour_data = 24'b110101111010100001001100;
		12'b011000100101: colour_data = 24'b110101111010100001001100;
		12'b011000100110: colour_data = 24'b110101111010100001001100;
		12'b011000100111: colour_data = 24'b110101111010100001001100;
		12'b011000101000: colour_data = 24'b110101111010100001001100;
		12'b011000101001: colour_data = 24'b110101111010100001001100;
		12'b011000101010: colour_data = 24'b110101111010100001001100;
		12'b011000101011: colour_data = 24'b110101111010100001001100;
		12'b011000101100: colour_data = 24'b110101111010100001001100;
		12'b011000101101: colour_data = 24'b110101111010100001001100;
		12'b011000101110: colour_data = 24'b110101111010100001001100;
		12'b011000101111: colour_data = 24'b110101111010100001001100;
		12'b011000110000: colour_data = 24'b110101111010100001001100;
		12'b011000110001: colour_data = 24'b110101111010100001001100;
		12'b011000110010: colour_data = 24'b110101111010100001001100;
		12'b011000110011: colour_data = 24'b110101111010100001001100;
		12'b011000110100: colour_data = 24'b110101111010100001001100;
		12'b011000110101: colour_data = 24'b110101111010100001001100;
		12'b011000110110: colour_data = 24'b110101111010100001001100;
		12'b011000110111: colour_data = 24'b110101111010100001001100;
		12'b011000111000: colour_data = 24'b110101111010100001001100;
		12'b011000111001: colour_data = 24'b110101111010100001001100;
		12'b011000111010: colour_data = 24'b110101111010100001001100;
		12'b011000111011: colour_data = 24'b110101111010100001001100;
		12'b011000111100: colour_data = 24'b110101111010100001001100;
		12'b011000111101: colour_data = 24'b110101111010100001001100;
		12'b011000111110: colour_data = 24'b110101111010100001001100;
		12'b011000111111: colour_data = 24'b110101111010100001001100;
		12'b011001000000: colour_data = 24'b110101111010100001001100;
		12'b011001000001: colour_data = 24'b110101111010100001001100;
		12'b011001000010: colour_data = 24'b110101111010100001001100;
		12'b011001000011: colour_data = 24'b110101111010100001001100;
		12'b011001000100: colour_data = 24'b110101111010100001001100;
		12'b011001000101: colour_data = 24'b110101111010100001001100;
		12'b011001000110: colour_data = 24'b110101111010100001001100;
		12'b011001000111: colour_data = 24'b110101111010100001001100;
		12'b011001001000: colour_data = 24'b110101111010100001001100;
		12'b011001001001: colour_data = 24'b110101111010100001001100;
		12'b011001001010: colour_data = 24'b110101111010100001001100;
		12'b011001001011: colour_data = 24'b110101111010100001001100;
		12'b011001001100: colour_data = 24'b110101111010100001001100;
		12'b011001001101: colour_data = 24'b110101111010100001001100;
		12'b011001001110: colour_data = 24'b110101111010100001001100;
		12'b011001001111: colour_data = 24'b110101111010100001001100;
		12'b011001010000: colour_data = 24'b110101111010100001001100;
		12'b011001010001: colour_data = 24'b110101111010100001001100;
		12'b011001010010: colour_data = 24'b110101111010100001001100;
		12'b011001010011: colour_data = 24'b110101111010100001001100;
		12'b011001010100: colour_data = 24'b110101111010100001001100;
		12'b011001010101: colour_data = 24'b110101111010100001001100;
		12'b011001010110: colour_data = 24'b110101111010100001001100;
		12'b011001010111: colour_data = 24'b110101111010100001001100;
		12'b011001011000: colour_data = 24'b110101111010100001001100;
		12'b011001011001: colour_data = 24'b110101111010100001001100;
		12'b011001011010: colour_data = 24'b110101111010100001001100;
		12'b011001011011: colour_data = 24'b110101111010100001001100;
		12'b011001011100: colour_data = 24'b110101111010100001001100;
		12'b011001011101: colour_data = 24'b110101111010100001001100;
		12'b011001011110: colour_data = 24'b110101111010100001001100;
		12'b011001011111: colour_data = 24'b110101111010100001001100;
		12'b011001100000: colour_data = 24'b110101111010100001001100;
		12'b011001100001: colour_data = 24'b110101111010100001001100;
		12'b011001100010: colour_data = 24'b110101111010100001001100;
		12'b011001100011: colour_data = 24'b110101111010100001001100;
		12'b011001100100: colour_data = 24'b110101111010100001001100;
		12'b011001100101: colour_data = 24'b110101111010100001001100;
		12'b011001100110: colour_data = 24'b110101111010100001001100;
		12'b011001100111: colour_data = 24'b110101111010100001001100;
		12'b011001101000: colour_data = 24'b110101111010100001001100;
		12'b011001101001: colour_data = 24'b110101111010100001001100;
		12'b011001101010: colour_data = 24'b110101111010100001001100;
		12'b011001101011: colour_data = 24'b110101111010100001001100;
		12'b011001101100: colour_data = 24'b110101111010100001001100;
		12'b011001101101: colour_data = 24'b110101111010100001001100;
		12'b011001101110: colour_data = 24'b110101111010100001001100;
		12'b011001101111: colour_data = 24'b110101111010100001001100;
		12'b011001110000: colour_data = 24'b110101111010100001001100;
		12'b011001110001: colour_data = 24'b110101111010100001001100;
		12'b011001110010: colour_data = 24'b110101111010100001001100;
		12'b011001110011: colour_data = 24'b110101111010100001001100;
		12'b011001110100: colour_data = 24'b110101111010100001001100;
		12'b011001110101: colour_data = 24'b110101111010100001001100;
		12'b011001110110: colour_data = 24'b110101111010100001001100;
		12'b011001110111: colour_data = 24'b110101111010100001001100;
		12'b011001111000: colour_data = 24'b110101111010100001001100;
		12'b011001111001: colour_data = 24'b110101111010100001001100;
		12'b011001111010: colour_data = 24'b110101111010100001001100;
		12'b011001111011: colour_data = 24'b110101111010100001001100;
		12'b011001111100: colour_data = 24'b110101111010100001001100;
		12'b011001111101: colour_data = 24'b110101111010100001001100;
		12'b011001111110: colour_data = 24'b110101111010100001001100;
		12'b011001111111: colour_data = 24'b110101111010100001001100;
		12'b011010000000: colour_data = 24'b110101111010100001001100;
		12'b011010000001: colour_data = 24'b110101111010100001001100;
		12'b011010000010: colour_data = 24'b110101111010100001001100;
		12'b011010000011: colour_data = 24'b110101111010100001001100;
		12'b011010000100: colour_data = 24'b110101111010100001001100;
		12'b011010000101: colour_data = 24'b110101111010100001001100;
		12'b011010000110: colour_data = 24'b110101111010100001001100;
		12'b011010000111: colour_data = 24'b110101111010100001001100;
		12'b011010001000: colour_data = 24'b110101111010100001001100;
		12'b011010001001: colour_data = 24'b110101111010100001001100;
		12'b011010001010: colour_data = 24'b110101111010100001001100;
		12'b011010001011: colour_data = 24'b110101111010100001001100;

		12'b011100000000: colour_data = 24'b110111101101100010010101;
		12'b011100000001: colour_data = 24'b110111101101100010010101;
		12'b011100000010: colour_data = 24'b110111101101100010010101;
		12'b011100000011: colour_data = 24'b110111101101100010010101;
		12'b011100000100: colour_data = 24'b110111101101100010010101;
		12'b011100000101: colour_data = 24'b110111101101100010010101;
		12'b011100000110: colour_data = 24'b110111101101100010010101;
		12'b011100000111: colour_data = 24'b110111101101100010010101;
		12'b011100001000: colour_data = 24'b110111101101100010010101;
		12'b011100001001: colour_data = 24'b110111101101100010010101;
		12'b011100001010: colour_data = 24'b110111101101100010010101;
		12'b011100001011: colour_data = 24'b110111101101100010010101;
		12'b011100001100: colour_data = 24'b110111101101100010010101;
		12'b011100001101: colour_data = 24'b110111101101100010010101;
		12'b011100001110: colour_data = 24'b110111101101100010010101;
		12'b011100001111: colour_data = 24'b110111101101100010010101;
		12'b011100010000: colour_data = 24'b110111101101100010010101;
		12'b011100010001: colour_data = 24'b110111101101100010010101;
		12'b011100010010: colour_data = 24'b110111101101100010010101;
		12'b011100010011: colour_data = 24'b110111101101100010010101;
		12'b011100010100: colour_data = 24'b110111101101100010010101;
		12'b011100010101: colour_data = 24'b110111101101100010010101;
		12'b011100010110: colour_data = 24'b110111101101100010010101;
		12'b011100010111: colour_data = 24'b110111101101100010010101;
		12'b011100011000: colour_data = 24'b110111101101100010010101;
		12'b011100011001: colour_data = 24'b110111101101100010010101;
		12'b011100011010: colour_data = 24'b110111101101100010010101;
		12'b011100011011: colour_data = 24'b110111101101100010010101;
		12'b011100011100: colour_data = 24'b110111101101100010010101;
		12'b011100011101: colour_data = 24'b110111101101100010010101;
		12'b011100011110: colour_data = 24'b110111101101100010010101;
		12'b011100011111: colour_data = 24'b110111101101100010010101;
		12'b011100100000: colour_data = 24'b110111101101100010010101;
		12'b011100100001: colour_data = 24'b110111101101100010010101;
		12'b011100100010: colour_data = 24'b110111101101100010010101;
		12'b011100100011: colour_data = 24'b110111101101100010010101;
		12'b011100100100: colour_data = 24'b110111101101100010010101;
		12'b011100100101: colour_data = 24'b110111101101100010010101;
		12'b011100100110: colour_data = 24'b110111101101100010010101;
		12'b011100100111: colour_data = 24'b110111101101100010010101;
		12'b011100101000: colour_data = 24'b110111101101100010010101;
		12'b011100101001: colour_data = 24'b110111101101100010010101;
		12'b011100101010: colour_data = 24'b110111101101100010010101;
		12'b011100101011: colour_data = 24'b110111101101100010010101;
		12'b011100101100: colour_data = 24'b110111101101100010010101;
		12'b011100101101: colour_data = 24'b110111101101100010010101;
		12'b011100101110: colour_data = 24'b110111101101100010010101;
		12'b011100101111: colour_data = 24'b110111101101100010010101;
		12'b011100110000: colour_data = 24'b110111101101100010010101;
		12'b011100110001: colour_data = 24'b110111101101100010010101;
		12'b011100110010: colour_data = 24'b110111101101100010010101;
		12'b011100110011: colour_data = 24'b110111101101100010010101;
		12'b011100110100: colour_data = 24'b110111101101100010010101;
		12'b011100110101: colour_data = 24'b110111101101100010010101;
		12'b011100110110: colour_data = 24'b110111101101100010010101;
		12'b011100110111: colour_data = 24'b110111101101100010010101;
		12'b011100111000: colour_data = 24'b110111101101100010010101;
		12'b011100111001: colour_data = 24'b110111101101100010010101;
		12'b011100111010: colour_data = 24'b110111101101100010010101;
		12'b011100111011: colour_data = 24'b110111101101100010010101;
		12'b011100111100: colour_data = 24'b110111101101100010010101;
		12'b011100111101: colour_data = 24'b110111101101100010010101;
		12'b011100111110: colour_data = 24'b110111101101100010010101;
		12'b011100111111: colour_data = 24'b110111101101100010010101;
		12'b011101000000: colour_data = 24'b110111101101100010010101;
		12'b011101000001: colour_data = 24'b110111101101100010010101;
		12'b011101000010: colour_data = 24'b110111101101100010010101;
		12'b011101000011: colour_data = 24'b110111101101100010010101;
		12'b011101000100: colour_data = 24'b110111101101100010010101;
		12'b011101000101: colour_data = 24'b110111101101100010010101;
		12'b011101000110: colour_data = 24'b110111101101100010010101;
		12'b011101000111: colour_data = 24'b110111101101100010010101;
		12'b011101001000: colour_data = 24'b110111101101100010010101;
		12'b011101001001: colour_data = 24'b110111101101100010010101;
		12'b011101001010: colour_data = 24'b110111101101100010010101;
		12'b011101001011: colour_data = 24'b110111101101100010010101;
		12'b011101001100: colour_data = 24'b110111101101100010010101;
		12'b011101001101: colour_data = 24'b110111101101100010010101;
		12'b011101001110: colour_data = 24'b110111101101100010010101;
		12'b011101001111: colour_data = 24'b110111101101100010010101;
		12'b011101010000: colour_data = 24'b110111101101100010010101;
		12'b011101010001: colour_data = 24'b110111101101100010010101;
		12'b011101010010: colour_data = 24'b110111101101100010010101;
		12'b011101010011: colour_data = 24'b110111101101100010010101;
		12'b011101010100: colour_data = 24'b110111101101100010010101;
		12'b011101010101: colour_data = 24'b110111101101100010010101;
		12'b011101010110: colour_data = 24'b110111101101100010010101;
		12'b011101010111: colour_data = 24'b110111101101100010010101;
		12'b011101011000: colour_data = 24'b110111101101100010010101;
		12'b011101011001: colour_data = 24'b110111101101100010010101;
		12'b011101011010: colour_data = 24'b110111101101100010010101;
		12'b011101011011: colour_data = 24'b110111101101100010010101;
		12'b011101011100: colour_data = 24'b110111101101100010010101;
		12'b011101011101: colour_data = 24'b110111101101100010010101;
		12'b011101011110: colour_data = 24'b110111101101100010010101;
		12'b011101011111: colour_data = 24'b110111101101100010010101;
		12'b011101100000: colour_data = 24'b110111101101100010010101;
		12'b011101100001: colour_data = 24'b110111101101100010010101;
		12'b011101100010: colour_data = 24'b110111101101100010010101;
		12'b011101100011: colour_data = 24'b110111101101100010010101;
		12'b011101100100: colour_data = 24'b110111101101100010010101;
		12'b011101100101: colour_data = 24'b110111101101100010010101;
		12'b011101100110: colour_data = 24'b110111101101100010010101;
		12'b011101100111: colour_data = 24'b110111101101100010010101;
		12'b011101101000: colour_data = 24'b110111101101100010010101;
		12'b011101101001: colour_data = 24'b110111101101100010010101;
		12'b011101101010: colour_data = 24'b110111101101100010010101;
		12'b011101101011: colour_data = 24'b110111101101100010010101;
		12'b011101101100: colour_data = 24'b110111101101100010010101;
		12'b011101101101: colour_data = 24'b110111101101100010010101;
		12'b011101101110: colour_data = 24'b110111101101100010010101;
		12'b011101101111: colour_data = 24'b110111101101100010010101;
		12'b011101110000: colour_data = 24'b110111101101100010010101;
		12'b011101110001: colour_data = 24'b110111101101100010010101;
		12'b011101110010: colour_data = 24'b110111101101100010010101;
		12'b011101110011: colour_data = 24'b110111101101100010010101;
		12'b011101110100: colour_data = 24'b110111101101100010010101;
		12'b011101110101: colour_data = 24'b110111101101100010010101;
		12'b011101110110: colour_data = 24'b110111101101100010010101;
		12'b011101110111: colour_data = 24'b110111101101100010010101;
		12'b011101111000: colour_data = 24'b110111101101100010010101;
		12'b011101111001: colour_data = 24'b110111101101100010010101;
		12'b011101111010: colour_data = 24'b110111101101100010010101;
		12'b011101111011: colour_data = 24'b110111101101100010010101;
		12'b011101111100: colour_data = 24'b110111101101100010010101;
		12'b011101111101: colour_data = 24'b110111101101100010010101;
		12'b011101111110: colour_data = 24'b110111101101100010010101;
		12'b011101111111: colour_data = 24'b110111101101100010010101;
		12'b011110000000: colour_data = 24'b110111101101100010010101;
		12'b011110000001: colour_data = 24'b110111101101100010010101;
		12'b011110000010: colour_data = 24'b110111101101100010010101;
		12'b011110000011: colour_data = 24'b110111101101100010010101;
		12'b011110000100: colour_data = 24'b110111101101100010010101;
		12'b011110000101: colour_data = 24'b110111101101100010010101;
		12'b011110000110: colour_data = 24'b110111101101100010010101;
		12'b011110000111: colour_data = 24'b110111101101100010010101;
		12'b011110001000: colour_data = 24'b110111101101100010010101;
		12'b011110001001: colour_data = 24'b110111101101100010010101;
		12'b011110001010: colour_data = 24'b110111101101100010010101;
		12'b011110001011: colour_data = 24'b110111101101100010010101;

		12'b100000000000: colour_data = 24'b110111101101100010010101;
		12'b100000000001: colour_data = 24'b110111101101100010010101;
		12'b100000000010: colour_data = 24'b110111101101100010010101;
		12'b100000000011: colour_data = 24'b110111101101100010010101;
		12'b100000000100: colour_data = 24'b110111101101100010010101;
		12'b100000000101: colour_data = 24'b110111101101100010010101;
		12'b100000000110: colour_data = 24'b110111101101100010010101;
		12'b100000000111: colour_data = 24'b110111101101100010010101;
		12'b100000001000: colour_data = 24'b110111101101100010010101;
		12'b100000001001: colour_data = 24'b110111101101100010010101;
		12'b100000001010: colour_data = 24'b110111101101100010010101;
		12'b100000001011: colour_data = 24'b110111101101100010010101;
		12'b100000001100: colour_data = 24'b110111101101100010010101;
		12'b100000001101: colour_data = 24'b110111101101100010010101;
		12'b100000001110: colour_data = 24'b110111101101100010010101;
		12'b100000001111: colour_data = 24'b110111101101100010010101;
		12'b100000010000: colour_data = 24'b110111101101100010010101;
		12'b100000010001: colour_data = 24'b110111101101100010010101;
		12'b100000010010: colour_data = 24'b110111101101100010010101;
		12'b100000010011: colour_data = 24'b110111101101100010010101;
		12'b100000010100: colour_data = 24'b110111101101100010010101;
		12'b100000010101: colour_data = 24'b110111101101100010010101;
		12'b100000010110: colour_data = 24'b110111101101100010010101;
		12'b100000010111: colour_data = 24'b110111101101100010010101;
		12'b100000011000: colour_data = 24'b110111101101100010010101;
		12'b100000011001: colour_data = 24'b110111101101100010010101;
		12'b100000011010: colour_data = 24'b110111101101100010010101;
		12'b100000011011: colour_data = 24'b110111101101100010010101;
		12'b100000011100: colour_data = 24'b110111101101100010010101;
		12'b100000011101: colour_data = 24'b110111101101100010010101;
		12'b100000011110: colour_data = 24'b110111101101100010010101;
		12'b100000011111: colour_data = 24'b110111101101100010010101;
		12'b100000100000: colour_data = 24'b110111101101100010010101;
		12'b100000100001: colour_data = 24'b110111101101100010010101;
		12'b100000100010: colour_data = 24'b110111101101100010010101;
		12'b100000100011: colour_data = 24'b110111101101100010010101;
		12'b100000100100: colour_data = 24'b110111101101100010010101;
		12'b100000100101: colour_data = 24'b110111101101100010010101;
		12'b100000100110: colour_data = 24'b110111101101100010010101;
		12'b100000100111: colour_data = 24'b110111101101100010010101;
		12'b100000101000: colour_data = 24'b110111101101100010010101;
		12'b100000101001: colour_data = 24'b110111101101100010010101;
		12'b100000101010: colour_data = 24'b110111101101100010010101;
		12'b100000101011: colour_data = 24'b110111101101100010010101;
		12'b100000101100: colour_data = 24'b110111101101100010010101;
		12'b100000101101: colour_data = 24'b110111101101100010010101;
		12'b100000101110: colour_data = 24'b110111101101100010010101;
		12'b100000101111: colour_data = 24'b110111101101100010010101;
		12'b100000110000: colour_data = 24'b110111101101100010010101;
		12'b100000110001: colour_data = 24'b110111101101100010010101;
		12'b100000110010: colour_data = 24'b110111101101100010010101;
		12'b100000110011: colour_data = 24'b110111101101100010010101;
		12'b100000110100: colour_data = 24'b110111101101100010010101;
		12'b100000110101: colour_data = 24'b110111101101100010010101;
		12'b100000110110: colour_data = 24'b110111101101100010010101;
		12'b100000110111: colour_data = 24'b110111101101100010010101;
		12'b100000111000: colour_data = 24'b110111101101100010010101;
		12'b100000111001: colour_data = 24'b110111101101100010010101;
		12'b100000111010: colour_data = 24'b110111101101100010010101;
		12'b100000111011: colour_data = 24'b110111101101100010010101;
		12'b100000111100: colour_data = 24'b110111101101100010010101;
		12'b100000111101: colour_data = 24'b110111101101100010010101;
		12'b100000111110: colour_data = 24'b110111101101100010010101;
		12'b100000111111: colour_data = 24'b110111101101100010010101;
		12'b100001000000: colour_data = 24'b110111101101100010010101;
		12'b100001000001: colour_data = 24'b110111101101100010010101;
		12'b100001000010: colour_data = 24'b110111101101100010010101;
		12'b100001000011: colour_data = 24'b110111101101100010010101;
		12'b100001000100: colour_data = 24'b110111101101100010010101;
		12'b100001000101: colour_data = 24'b110111101101100010010101;
		12'b100001000110: colour_data = 24'b110111101101100010010101;
		12'b100001000111: colour_data = 24'b110111101101100010010101;
		12'b100001001000: colour_data = 24'b110111101101100010010101;
		12'b100001001001: colour_data = 24'b110111101101100010010101;
		12'b100001001010: colour_data = 24'b110111101101100010010101;
		12'b100001001011: colour_data = 24'b110111101101100010010101;
		12'b100001001100: colour_data = 24'b110111101101100010010101;
		12'b100001001101: colour_data = 24'b110111101101100010010101;
		12'b100001001110: colour_data = 24'b110111101101100010010101;
		12'b100001001111: colour_data = 24'b110111101101100010010101;
		12'b100001010000: colour_data = 24'b110111101101100010010101;
		12'b100001010001: colour_data = 24'b110111101101100010010101;
		12'b100001010010: colour_data = 24'b110111101101100010010101;
		12'b100001010011: colour_data = 24'b110111101101100010010101;
		12'b100001010100: colour_data = 24'b110111101101100010010101;
		12'b100001010101: colour_data = 24'b110111101101100010010101;
		12'b100001010110: colour_data = 24'b110111101101100010010101;
		12'b100001010111: colour_data = 24'b110111101101100010010101;
		12'b100001011000: colour_data = 24'b110111101101100010010101;
		12'b100001011001: colour_data = 24'b110111101101100010010101;
		12'b100001011010: colour_data = 24'b110111101101100010010101;
		12'b100001011011: colour_data = 24'b110111101101100010010101;
		12'b100001011100: colour_data = 24'b110111101101100010010101;
		12'b100001011101: colour_data = 24'b110111101101100010010101;
		12'b100001011110: colour_data = 24'b110111101101100010010101;
		12'b100001011111: colour_data = 24'b110111101101100010010101;
		12'b100001100000: colour_data = 24'b110111101101100010010101;
		12'b100001100001: colour_data = 24'b110111101101100010010101;
		12'b100001100010: colour_data = 24'b110111101101100010010101;
		12'b100001100011: colour_data = 24'b110111101101100010010101;
		12'b100001100100: colour_data = 24'b110111101101100010010101;
		12'b100001100101: colour_data = 24'b110111101101100010010101;
		12'b100001100110: colour_data = 24'b110111101101100010010101;
		12'b100001100111: colour_data = 24'b110111101101100010010101;
		12'b100001101000: colour_data = 24'b110111101101100010010101;
		12'b100001101001: colour_data = 24'b110111101101100010010101;
		12'b100001101010: colour_data = 24'b110111101101100010010101;
		12'b100001101011: colour_data = 24'b110111101101100010010101;
		12'b100001101100: colour_data = 24'b110111101101100010010101;
		12'b100001101101: colour_data = 24'b110111101101100010010101;
		12'b100001101110: colour_data = 24'b110111101101100010010101;
		12'b100001101111: colour_data = 24'b110111101101100010010101;
		12'b100001110000: colour_data = 24'b110111101101100010010101;
		12'b100001110001: colour_data = 24'b110111101101100010010101;
		12'b100001110010: colour_data = 24'b110111101101100010010101;
		12'b100001110011: colour_data = 24'b110111101101100010010101;
		12'b100001110100: colour_data = 24'b110111101101100010010101;
		12'b100001110101: colour_data = 24'b110111101101100010010101;
		12'b100001110110: colour_data = 24'b110111101101100010010101;
		12'b100001110111: colour_data = 24'b110111101101100010010101;
		12'b100001111000: colour_data = 24'b110111101101100010010101;
		12'b100001111001: colour_data = 24'b110111101101100010010101;
		12'b100001111010: colour_data = 24'b110111101101100010010101;
		12'b100001111011: colour_data = 24'b110111101101100010010101;
		12'b100001111100: colour_data = 24'b110111101101100010010101;
		12'b100001111101: colour_data = 24'b110111101101100010010101;
		12'b100001111110: colour_data = 24'b110111101101100010010101;
		12'b100001111111: colour_data = 24'b110111101101100010010101;
		12'b100010000000: colour_data = 24'b110111101101100010010101;
		12'b100010000001: colour_data = 24'b110111101101100010010101;
		12'b100010000010: colour_data = 24'b110111101101100010010101;
		12'b100010000011: colour_data = 24'b110111101101100010010101;
		12'b100010000100: colour_data = 24'b110111101101100010010101;
		12'b100010000101: colour_data = 24'b110111101101100010010101;
		12'b100010000110: colour_data = 24'b110111101101100010010101;
		12'b100010000111: colour_data = 24'b110111101101100010010101;
		12'b100010001000: colour_data = 24'b110111101101100010010101;
		12'b100010001001: colour_data = 24'b110111101101100010010101;
		12'b100010001010: colour_data = 24'b110111101101100010010101;
		12'b100010001011: colour_data = 24'b110111101101100010010101;

		12'b100100000000: colour_data = 24'b110111101101100010010101;
		12'b100100000001: colour_data = 24'b110111101101100010010101;
		12'b100100000010: colour_data = 24'b110111101101100010010101;
		12'b100100000011: colour_data = 24'b110111101101100010010101;
		12'b100100000100: colour_data = 24'b110111101101100010010101;
		12'b100100000101: colour_data = 24'b110111101101100010010101;
		12'b100100000110: colour_data = 24'b110111101101100010010101;
		12'b100100000111: colour_data = 24'b110111101101100010010101;
		12'b100100001000: colour_data = 24'b110111101101100010010101;
		12'b100100001001: colour_data = 24'b110111101101100010010101;
		12'b100100001010: colour_data = 24'b110111101101100010010101;
		12'b100100001011: colour_data = 24'b110111101101100010010101;
		12'b100100001100: colour_data = 24'b110111101101100010010101;
		12'b100100001101: colour_data = 24'b110111101101100010010101;
		12'b100100001110: colour_data = 24'b110111101101100010010101;
		12'b100100001111: colour_data = 24'b110111101101100010010101;
		12'b100100010000: colour_data = 24'b110111101101100010010101;
		12'b100100010001: colour_data = 24'b110111101101100010010101;
		12'b100100010010: colour_data = 24'b110111101101100010010101;
		12'b100100010011: colour_data = 24'b110111101101100010010101;
		12'b100100010100: colour_data = 24'b110111101101100010010101;
		12'b100100010101: colour_data = 24'b110111101101100010010101;
		12'b100100010110: colour_data = 24'b110111101101100010010101;
		12'b100100010111: colour_data = 24'b110111101101100010010101;
		12'b100100011000: colour_data = 24'b110111101101100010010101;
		12'b100100011001: colour_data = 24'b110111101101100010010101;
		12'b100100011010: colour_data = 24'b110111101101100010010101;
		12'b100100011011: colour_data = 24'b110111101101100010010101;
		12'b100100011100: colour_data = 24'b110111101101100010010101;
		12'b100100011101: colour_data = 24'b110111101101100010010101;
		12'b100100011110: colour_data = 24'b110111101101100010010101;
		12'b100100011111: colour_data = 24'b110111101101100010010101;
		12'b100100100000: colour_data = 24'b110111101101100010010101;
		12'b100100100001: colour_data = 24'b110111101101100010010101;
		12'b100100100010: colour_data = 24'b110111101101100010010101;
		12'b100100100011: colour_data = 24'b110111101101100010010101;
		12'b100100100100: colour_data = 24'b110111101101100010010101;
		12'b100100100101: colour_data = 24'b110111101101100010010101;
		12'b100100100110: colour_data = 24'b110111101101100010010101;
		12'b100100100111: colour_data = 24'b110111101101100010010101;
		12'b100100101000: colour_data = 24'b110111101101100010010101;
		12'b100100101001: colour_data = 24'b110111101101100010010101;
		12'b100100101010: colour_data = 24'b110111101101100010010101;
		12'b100100101011: colour_data = 24'b110111101101100010010101;
		12'b100100101100: colour_data = 24'b110111101101100010010101;
		12'b100100101101: colour_data = 24'b110111101101100010010101;
		12'b100100101110: colour_data = 24'b110111101101100010010101;
		12'b100100101111: colour_data = 24'b110111101101100010010101;
		12'b100100110000: colour_data = 24'b110111101101100010010101;
		12'b100100110001: colour_data = 24'b110111101101100010010101;
		12'b100100110010: colour_data = 24'b110111101101100010010101;
		12'b100100110011: colour_data = 24'b110111101101100010010101;
		12'b100100110100: colour_data = 24'b110111101101100010010101;
		12'b100100110101: colour_data = 24'b110111101101100010010101;
		12'b100100110110: colour_data = 24'b110111101101100010010101;
		12'b100100110111: colour_data = 24'b110111101101100010010101;
		12'b100100111000: colour_data = 24'b110111101101100010010101;
		12'b100100111001: colour_data = 24'b110111101101100010010101;
		12'b100100111010: colour_data = 24'b110111101101100010010101;
		12'b100100111011: colour_data = 24'b110111101101100010010101;
		12'b100100111100: colour_data = 24'b110111101101100010010101;
		12'b100100111101: colour_data = 24'b110111101101100010010101;
		12'b100100111110: colour_data = 24'b110111101101100010010101;
		12'b100100111111: colour_data = 24'b110111101101100010010101;
		12'b100101000000: colour_data = 24'b110111101101100010010101;
		12'b100101000001: colour_data = 24'b110111101101100010010101;
		12'b100101000010: colour_data = 24'b110111101101100010010101;
		12'b100101000011: colour_data = 24'b110111101101100010010101;
		12'b100101000100: colour_data = 24'b110111101101100010010101;
		12'b100101000101: colour_data = 24'b110111101101100010010101;
		12'b100101000110: colour_data = 24'b110111101101100010010101;
		12'b100101000111: colour_data = 24'b110111101101100010010101;
		12'b100101001000: colour_data = 24'b110111101101100010010101;
		12'b100101001001: colour_data = 24'b110111101101100010010101;
		12'b100101001010: colour_data = 24'b110111101101100010010101;
		12'b100101001011: colour_data = 24'b110111101101100010010101;
		12'b100101001100: colour_data = 24'b110111101101100010010101;
		12'b100101001101: colour_data = 24'b110111101101100010010101;
		12'b100101001110: colour_data = 24'b110111101101100010010101;
		12'b100101001111: colour_data = 24'b110111101101100010010101;
		12'b100101010000: colour_data = 24'b110111101101100010010101;
		12'b100101010001: colour_data = 24'b110111101101100010010101;
		12'b100101010010: colour_data = 24'b110111101101100010010101;
		12'b100101010011: colour_data = 24'b110111101101100010010101;
		12'b100101010100: colour_data = 24'b110111101101100010010101;
		12'b100101010101: colour_data = 24'b110111101101100010010101;
		12'b100101010110: colour_data = 24'b110111101101100010010101;
		12'b100101010111: colour_data = 24'b110111101101100010010101;
		12'b100101011000: colour_data = 24'b110111101101100010010101;
		12'b100101011001: colour_data = 24'b110111101101100010010101;
		12'b100101011010: colour_data = 24'b110111101101100010010101;
		12'b100101011011: colour_data = 24'b110111101101100010010101;
		12'b100101011100: colour_data = 24'b110111101101100010010101;
		12'b100101011101: colour_data = 24'b110111101101100010010101;
		12'b100101011110: colour_data = 24'b110111101101100010010101;
		12'b100101011111: colour_data = 24'b110111101101100010010101;
		12'b100101100000: colour_data = 24'b110111101101100010010101;
		12'b100101100001: colour_data = 24'b110111101101100010010101;
		12'b100101100010: colour_data = 24'b110111101101100010010101;
		12'b100101100011: colour_data = 24'b110111101101100010010101;
		12'b100101100100: colour_data = 24'b110111101101100010010101;
		12'b100101100101: colour_data = 24'b110111101101100010010101;
		12'b100101100110: colour_data = 24'b110111101101100010010101;
		12'b100101100111: colour_data = 24'b110111101101100010010101;
		12'b100101101000: colour_data = 24'b110111101101100010010101;
		12'b100101101001: colour_data = 24'b110111101101100010010101;
		12'b100101101010: colour_data = 24'b110111101101100010010101;
		12'b100101101011: colour_data = 24'b110111101101100010010101;
		12'b100101101100: colour_data = 24'b110111101101100010010101;
		12'b100101101101: colour_data = 24'b110111101101100010010101;
		12'b100101101110: colour_data = 24'b110111101101100010010101;
		12'b100101101111: colour_data = 24'b110111101101100010010101;
		12'b100101110000: colour_data = 24'b110111101101100010010101;
		12'b100101110001: colour_data = 24'b110111101101100010010101;
		12'b100101110010: colour_data = 24'b110111101101100010010101;
		12'b100101110011: colour_data = 24'b110111101101100010010101;
		12'b100101110100: colour_data = 24'b110111101101100010010101;
		12'b100101110101: colour_data = 24'b110111101101100010010101;
		12'b100101110110: colour_data = 24'b110111101101100010010101;
		12'b100101110111: colour_data = 24'b110111101101100010010101;
		12'b100101111000: colour_data = 24'b110111101101100010010101;
		12'b100101111001: colour_data = 24'b110111101101100010010101;
		12'b100101111010: colour_data = 24'b110111101101100010010101;
		12'b100101111011: colour_data = 24'b110111101101100010010101;
		12'b100101111100: colour_data = 24'b110111101101100010010101;
		12'b100101111101: colour_data = 24'b110111101101100010010101;
		12'b100101111110: colour_data = 24'b110111101101100010010101;
		12'b100101111111: colour_data = 24'b110111101101100010010101;
		12'b100110000000: colour_data = 24'b110111101101100010010101;
		12'b100110000001: colour_data = 24'b110111101101100010010101;
		12'b100110000010: colour_data = 24'b110111101101100010010101;
		12'b100110000011: colour_data = 24'b110111101101100010010101;
		12'b100110000100: colour_data = 24'b110111101101100010010101;
		12'b100110000101: colour_data = 24'b110111101101100010010101;
		12'b100110000110: colour_data = 24'b110111101101100010010101;
		12'b100110000111: colour_data = 24'b110111101101100010010101;
		12'b100110001000: colour_data = 24'b110111101101100010010101;
		12'b100110001001: colour_data = 24'b110111101101100010010101;
		12'b100110001010: colour_data = 24'b110111101101100010010101;
		12'b100110001011: colour_data = 24'b110111101101100010010101;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule