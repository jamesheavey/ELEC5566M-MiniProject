module character_physics#(
	parameter PLAYER_SIZE_X,
	parameter PLAYER_SIZE_Y
)(
	input GAME_clk, rst, flap,
	output reg [15:0] playerY,
	output reg [3:0] player_state
);

integer X_acc=2, Y_acc=2, X_vel_max=10, Y_vel_min=-20;
reg signed [15:0] X_vel, Y_vel;

always @(posedge GAME_clk or posedge rst)
begin
	if (rst) begin
		Y_vel <= 0;
		playerY <= (480 - PLAYER_SIZE_Y)/2;
	end else begin
		
		playerY <= playerY + Y_vel;
		
	end
end

endmodule
		