module sonic_run_2_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: colour_data = 24'b111111110000000010010110;
		12'b000000000001: colour_data = 24'b111111110000000010010110;
		12'b000000000010: colour_data = 24'b111111110000000010010110;
		12'b000000000011: colour_data = 24'b111111110000000010010110;
		12'b000000000100: colour_data = 24'b111111110000000010010110;
		12'b000000000101: colour_data = 24'b111111110000000010010110;
		12'b000000000110: colour_data = 24'b111111110000000010010110;
		12'b000000000111: colour_data = 24'b111111110000000010010110;
		12'b000000001000: colour_data = 24'b111111110000000010010110;
		12'b000000001001: colour_data = 24'b111111110000000010010110;
		12'b000000001010: colour_data = 24'b111111110000000010010110;
		12'b000000001011: colour_data = 24'b111111110000000010010110;
		12'b000000001100: colour_data = 24'b111111110000000010010110;
		12'b000000001101: colour_data = 24'b111111110000000010010110;
		12'b000000001110: colour_data = 24'b111111110000000010010110;
		12'b000000001111: colour_data = 24'b111111110000000010010110;
		12'b000000010000: colour_data = 24'b111111110000000010010110;
		12'b000000010001: colour_data = 24'b111111110000000010010110;
		12'b000000010010: colour_data = 24'b111111110000000010010110;
		12'b000000010011: colour_data = 24'b111111110000000010010110;
		12'b000000010100: colour_data = 24'b111111110000000010010110;
		12'b000000010101: colour_data = 24'b111111110000000010010110;
		12'b000000010110: colour_data = 24'b111111110000000010010110;
		12'b000000010111: colour_data = 24'b111111110000000010010110;
		12'b000000011000: colour_data = 24'b111111110000000010010110;
		12'b000000011001: colour_data = 24'b111111110000000010010110;
		12'b000000011010: colour_data = 24'b111111110000000010010110;
		12'b000000011011: colour_data = 24'b111111110000000010010110;
		12'b000000011100: colour_data = 24'b111111110000000010010110;
		12'b000000011101: colour_data = 24'b111111110000000010010110;
		12'b000000011110: colour_data = 24'b111111110000000010010110;
		12'b000000011111: colour_data = 24'b111111110000000010010110;
		12'b000000100000: colour_data = 24'b111111110000000010010110;
		12'b000000100001: colour_data = 24'b111111110000000010010110;
		12'b000000100010: colour_data = 24'b111111110000000010010110;
		12'b000000100011: colour_data = 24'b111111110000000010010110;
		12'b000000100100: colour_data = 24'b111111110000000010010110;

		12'b000001000000: colour_data = 24'b111111110000000010010110;
		12'b000001000001: colour_data = 24'b111111110000000010010110;
		12'b000001000010: colour_data = 24'b111111110000000010010110;
		12'b000001000011: colour_data = 24'b111111110000000010010110;
		12'b000001000100: colour_data = 24'b111111110000000010010110;
		12'b000001000101: colour_data = 24'b111111110000000010010110;
		12'b000001000110: colour_data = 24'b111111110000000010010110;
		12'b000001000111: colour_data = 24'b111111110000000010010110;
		12'b000001001000: colour_data = 24'b111111110000000010010110;
		12'b000001001001: colour_data = 24'b111111110000000010010110;
		12'b000001001010: colour_data = 24'b111111110000000010010110;
		12'b000001001011: colour_data = 24'b111111110000000010010110;
		12'b000001001100: colour_data = 24'b111111110000000010010110;
		12'b000001001101: colour_data = 24'b111111110000000010010110;
		12'b000001001110: colour_data = 24'b111111110000000010010110;
		12'b000001001111: colour_data = 24'b111111110000000010010110;
		12'b000001010000: colour_data = 24'b111111110000000010010110;
		12'b000001010001: colour_data = 24'b111111110000000010010110;
		12'b000001010010: colour_data = 24'b111111110000000010010110;
		12'b000001010011: colour_data = 24'b111111110000000010010110;
		12'b000001010100: colour_data = 24'b111111110000000010010110;
		12'b000001010101: colour_data = 24'b111111110000000010010110;
		12'b000001010110: colour_data = 24'b111111110000000010010110;
		12'b000001010111: colour_data = 24'b111111110000000010010110;
		12'b000001011000: colour_data = 24'b111111110000000010010110;
		12'b000001011001: colour_data = 24'b111111110000000010010110;
		12'b000001011010: colour_data = 24'b111111110000000010010110;
		12'b000001011011: colour_data = 24'b111111110000000010010110;
		12'b000001011100: colour_data = 24'b111111110000000010010110;
		12'b000001011101: colour_data = 24'b111111110000000010010110;
		12'b000001011110: colour_data = 24'b111111110000000010010110;
		12'b000001011111: colour_data = 24'b111111110000000010010110;
		12'b000001100000: colour_data = 24'b111111110000000010010110;
		12'b000001100001: colour_data = 24'b111111110000000010010110;
		12'b000001100010: colour_data = 24'b111111110000000010010110;
		12'b000001100011: colour_data = 24'b111111110000000010010110;
		12'b000001100100: colour_data = 24'b111111110000000010010110;

		12'b000010000000: colour_data = 24'b111111110000000010010110;
		12'b000010000001: colour_data = 24'b111111110000000010010110;
		12'b000010000010: colour_data = 24'b111111110000000010010110;
		12'b000010000011: colour_data = 24'b111111110000000010010110;
		12'b000010000100: colour_data = 24'b111111110000000010010110;
		12'b000010000101: colour_data = 24'b111111110000000010010110;
		12'b000010000110: colour_data = 24'b111111110000000010010110;
		12'b000010000111: colour_data = 24'b111111110000000010010110;
		12'b000010001000: colour_data = 24'b111111110000000010010110;
		12'b000010001001: colour_data = 24'b111111110000000010010110;
		12'b000010001010: colour_data = 24'b111111110000000010010110;
		12'b000010001011: colour_data = 24'b111111110000000010010110;
		12'b000010001100: colour_data = 24'b111111110000000010010110;
		12'b000010001101: colour_data = 24'b111111110000000010010110;
		12'b000010001110: colour_data = 24'b111111110000000010010110;
		12'b000010001111: colour_data = 24'b111111110000000010010110;
		12'b000010010000: colour_data = 24'b111111110000000010010110;
		12'b000010010001: colour_data = 24'b111111110000000010010110;
		12'b000010010010: colour_data = 24'b111111110000000010010110;
		12'b000010010011: colour_data = 24'b111111110000000010010110;
		12'b000010010100: colour_data = 24'b111111110000000010010110;
		12'b000010010101: colour_data = 24'b111111110000000010010110;
		12'b000010010110: colour_data = 24'b111111110000000010010110;
		12'b000010010111: colour_data = 24'b111111110000000010010110;
		12'b000010011000: colour_data = 24'b111111110000000010010110;
		12'b000010011001: colour_data = 24'b111111110000000010010110;
		12'b000010011010: colour_data = 24'b111111110000000010010110;
		12'b000010011011: colour_data = 24'b111111110000000010010110;
		12'b000010011100: colour_data = 24'b111111110000000010010110;
		12'b000010011101: colour_data = 24'b111111110000000010010110;
		12'b000010011110: colour_data = 24'b111111110000000010010110;
		12'b000010011111: colour_data = 24'b111111110000000010010110;
		12'b000010100000: colour_data = 24'b111111110000000010010110;
		12'b000010100001: colour_data = 24'b111111110000000010010110;
		12'b000010100010: colour_data = 24'b111111110000000010010110;
		12'b000010100011: colour_data = 24'b111111110000000010010110;
		12'b000010100100: colour_data = 24'b111111110000000010010110;

		12'b000011000000: colour_data = 24'b111111110000000010010110;
		12'b000011000001: colour_data = 24'b111111110000000010010110;
		12'b000011000010: colour_data = 24'b111111110000000010010110;
		12'b000011000011: colour_data = 24'b111111110000000010010110;
		12'b000011000100: colour_data = 24'b111111110000000010010110;
		12'b000011000101: colour_data = 24'b111111110000000010010110;
		12'b000011000110: colour_data = 24'b111111110000000010010110;
		12'b000011000111: colour_data = 24'b111111110000000010010110;
		12'b000011001000: colour_data = 24'b111111110000000010010110;
		12'b000011001001: colour_data = 24'b111111110000000010010110;
		12'b000011001010: colour_data = 24'b111111110000000010010110;
		12'b000011001011: colour_data = 24'b111111110000000010010110;
		12'b000011001100: colour_data = 24'b111111110000000010010110;
		12'b000011001101: colour_data = 24'b111111110000000010010110;
		12'b000011001110: colour_data = 24'b111111110000000010010110;
		12'b000011001111: colour_data = 24'b111111110000000010010110;
		12'b000011010000: colour_data = 24'b111111110000000010010110;
		12'b000011010001: colour_data = 24'b111111110000000010010110;
		12'b000011010010: colour_data = 24'b111111110000000010010110;
		12'b000011010011: colour_data = 24'b111111110000000010010110;
		12'b000011010100: colour_data = 24'b111111110000000010010110;
		12'b000011010101: colour_data = 24'b111111110000000010010110;
		12'b000011010110: colour_data = 24'b111111110000000010010110;
		12'b000011010111: colour_data = 24'b111111110000000010010110;
		12'b000011011000: colour_data = 24'b111111110000000010010110;
		12'b000011011001: colour_data = 24'b111111110000000010010110;
		12'b000011011010: colour_data = 24'b111111110000000010010110;
		12'b000011011011: colour_data = 24'b111111110000000010010110;
		12'b000011011100: colour_data = 24'b111111110000000010010110;
		12'b000011011101: colour_data = 24'b111111110000000010010110;
		12'b000011011110: colour_data = 24'b111111110000000010010110;
		12'b000011011111: colour_data = 24'b111111110000000010010110;
		12'b000011100000: colour_data = 24'b111111110000000010010110;
		12'b000011100001: colour_data = 24'b111111110000000010010110;
		12'b000011100010: colour_data = 24'b111111110000000010010110;
		12'b000011100011: colour_data = 24'b111111110000000010010110;
		12'b000011100100: colour_data = 24'b111111110000000010010110;

		12'b000100000000: colour_data = 24'b111111110000000010010110;
		12'b000100000001: colour_data = 24'b111111110000000010010110;
		12'b000100000010: colour_data = 24'b111111110000000010010110;
		12'b000100000011: colour_data = 24'b111111110000000010010110;
		12'b000100000100: colour_data = 24'b111111110000000010010110;
		12'b000100000101: colour_data = 24'b111111110000000010010110;
		12'b000100000110: colour_data = 24'b111111110000000010010110;
		12'b000100000111: colour_data = 24'b111111110000000010010110;
		12'b000100001000: colour_data = 24'b111111110000000010010110;
		12'b000100001001: colour_data = 24'b111111110000000010010110;
		12'b000100001010: colour_data = 24'b111111110000000010010110;
		12'b000100001011: colour_data = 24'b111111110000000010010110;
		12'b000100001100: colour_data = 24'b111111110000000010010110;
		12'b000100001101: colour_data = 24'b111111110000000010010110;
		12'b000100001110: colour_data = 24'b100010001000100011101110;
		12'b000100001111: colour_data = 24'b100010001000100011101110;
		12'b000100010000: colour_data = 24'b100010001000100011101110;
		12'b000100010001: colour_data = 24'b100010001000100011101110;
		12'b000100010010: colour_data = 24'b100010001000100011101110;
		12'b000100010011: colour_data = 24'b111111110000000010010110;
		12'b000100010100: colour_data = 24'b111111110000000010010110;
		12'b000100010101: colour_data = 24'b111111110000000010010110;
		12'b000100010110: colour_data = 24'b111111110000000010010110;
		12'b000100010111: colour_data = 24'b111111110000000010010110;
		12'b000100011000: colour_data = 24'b111111110000000010010110;
		12'b000100011001: colour_data = 24'b111111110000000010010110;
		12'b000100011010: colour_data = 24'b111111110000000010010110;
		12'b000100011011: colour_data = 24'b111111110000000010010110;
		12'b000100011100: colour_data = 24'b111111110000000010010110;
		12'b000100011101: colour_data = 24'b111111110000000010010110;
		12'b000100011110: colour_data = 24'b111111110000000010010110;
		12'b000100011111: colour_data = 24'b111111110000000010010110;
		12'b000100100000: colour_data = 24'b111111110000000010010110;
		12'b000100100001: colour_data = 24'b111111110000000010010110;
		12'b000100100010: colour_data = 24'b111111110000000010010110;
		12'b000100100011: colour_data = 24'b111111110000000010010110;
		12'b000100100100: colour_data = 24'b111111110000000010010110;

		12'b000101000000: colour_data = 24'b111111110000000010010110;
		12'b000101000001: colour_data = 24'b111111110000000010010110;
		12'b000101000010: colour_data = 24'b111111110000000010010110;
		12'b000101000011: colour_data = 24'b111111110000000010010110;
		12'b000101000100: colour_data = 24'b111111110000000010010110;
		12'b000101000101: colour_data = 24'b111111110000000010010110;
		12'b000101000110: colour_data = 24'b111111110000000010010110;
		12'b000101000111: colour_data = 24'b111111110000000010010110;
		12'b000101001000: colour_data = 24'b111111110000000010010110;
		12'b000101001001: colour_data = 24'b111111110000000010010110;
		12'b000101001010: colour_data = 24'b111111110000000010010110;
		12'b000101001011: colour_data = 24'b100010001000100011101110;
		12'b000101001100: colour_data = 24'b100010001000100011101110;
		12'b000101001101: colour_data = 24'b100010001000100011101110;
		12'b000101001110: colour_data = 24'b011001100110011011101110;
		12'b000101001111: colour_data = 24'b010001000100010011101110;
		12'b000101010000: colour_data = 24'b010001000100010011101110;
		12'b000101010001: colour_data = 24'b010001000100010011101110;
		12'b000101010010: colour_data = 24'b011001100110011011101110;
		12'b000101010011: colour_data = 24'b100010001000100011101110;
		12'b000101010100: colour_data = 24'b100010001000100011101110;
		12'b000101010101: colour_data = 24'b100010001000100011101110;
		12'b000101010110: colour_data = 24'b111111110000000010010110;
		12'b000101010111: colour_data = 24'b111111110000000010010110;
		12'b000101011000: colour_data = 24'b111111110000000010010110;
		12'b000101011001: colour_data = 24'b111111110000000010010110;
		12'b000101011010: colour_data = 24'b111111110000000010010110;
		12'b000101011011: colour_data = 24'b111111110000000010010110;
		12'b000101011100: colour_data = 24'b111111110000000010010110;
		12'b000101011101: colour_data = 24'b111111110000000010010110;
		12'b000101011110: colour_data = 24'b111111110000000010010110;
		12'b000101011111: colour_data = 24'b111111110000000010010110;
		12'b000101100000: colour_data = 24'b111111110000000010010110;
		12'b000101100001: colour_data = 24'b111111110000000010010110;
		12'b000101100010: colour_data = 24'b111111110000000010010110;
		12'b000101100011: colour_data = 24'b111111110000000010010110;
		12'b000101100100: colour_data = 24'b111111110000000010010110;

		12'b000110000000: colour_data = 24'b111111110000000010010110;
		12'b000110000001: colour_data = 24'b111111110000000010010110;
		12'b000110000010: colour_data = 24'b111111110000000010010110;
		12'b000110000011: colour_data = 24'b111111110000000010010110;
		12'b000110000100: colour_data = 24'b111111110000000010010110;
		12'b000110000101: colour_data = 24'b111111110000000010010110;
		12'b000110000110: colour_data = 24'b111111110000000010010110;
		12'b000110000111: colour_data = 24'b111111110000000010010110;
		12'b000110001000: colour_data = 24'b111111110000000010010110;
		12'b000110001001: colour_data = 24'b100010001000100011101110;
		12'b000110001010: colour_data = 24'b100010001000100011101110;
		12'b000110001011: colour_data = 24'b010001000100010011101110;
		12'b000110001100: colour_data = 24'b010001000100010011101110;
		12'b000110001101: colour_data = 24'b010001000100010011101110;
		12'b000110001110: colour_data = 24'b010001000100010011101110;
		12'b000110001111: colour_data = 24'b001000100010001011001100;
		12'b000110010000: colour_data = 24'b001000100010001011001100;
		12'b000110010001: colour_data = 24'b001000100010001011001100;
		12'b000110010010: colour_data = 24'b010001000100010011101110;
		12'b000110010011: colour_data = 24'b010001000100010011101110;
		12'b000110010100: colour_data = 24'b010001000100010011101110;
		12'b000110010101: colour_data = 24'b011001100110011011101110;
		12'b000110010110: colour_data = 24'b100010001000100011101110;
		12'b000110010111: colour_data = 24'b100010001000100011101110;
		12'b000110011000: colour_data = 24'b111111110000000010010110;
		12'b000110011001: colour_data = 24'b111111110000000010010110;
		12'b000110011010: colour_data = 24'b111111110000000010010110;
		12'b000110011011: colour_data = 24'b111111110000000010010110;
		12'b000110011100: colour_data = 24'b111111110000000010010110;
		12'b000110011101: colour_data = 24'b111111110000000010010110;
		12'b000110011110: colour_data = 24'b111111110000000010010110;
		12'b000110011111: colour_data = 24'b111111110000000010010110;
		12'b000110100000: colour_data = 24'b111111110000000010010110;
		12'b000110100001: colour_data = 24'b111111110000000010010110;
		12'b000110100010: colour_data = 24'b111111110000000010010110;
		12'b000110100011: colour_data = 24'b111111110000000010010110;
		12'b000110100100: colour_data = 24'b111111110000000010010110;

		12'b000111000000: colour_data = 24'b111111110000000010010110;
		12'b000111000001: colour_data = 24'b111111110000000010010110;
		12'b000111000010: colour_data = 24'b111111110000000010010110;
		12'b000111000011: colour_data = 24'b111111110000000010010110;
		12'b000111000100: colour_data = 24'b111111110000000010010110;
		12'b000111000101: colour_data = 24'b111111110000000010010110;
		12'b000111000110: colour_data = 24'b111111110000000010010110;
		12'b000111000111: colour_data = 24'b111111110000000010010110;
		12'b000111001000: colour_data = 24'b111111110000000010010110;
		12'b000111001001: colour_data = 24'b111111110000000010010110;
		12'b000111001010: colour_data = 24'b111111110000000010010110;
		12'b000111001011: colour_data = 24'b001000100010001011001100;
		12'b000111001100: colour_data = 24'b001000100010001011001100;
		12'b000111001101: colour_data = 24'b001000100010001011001100;
		12'b000111001110: colour_data = 24'b001000100010001011001100;
		12'b000111001111: colour_data = 24'b001000100010001011001100;
		12'b000111010000: colour_data = 24'b001000100010001011001100;
		12'b000111010001: colour_data = 24'b001000100010001011001100;
		12'b000111010010: colour_data = 24'b001000100010001011001100;
		12'b000111010011: colour_data = 24'b101101000110110001001000;
		12'b000111010100: colour_data = 24'b010001000100010011101110;
		12'b000111010101: colour_data = 24'b010001000100010011101110;
		12'b000111010110: colour_data = 24'b010001000100010011101110;
		12'b000111010111: colour_data = 24'b011001100110011011101110;
		12'b000111011000: colour_data = 24'b100010001000100011101110;
		12'b000111011001: colour_data = 24'b100010001000100011101110;
		12'b000111011010: colour_data = 24'b111111110000000010010110;
		12'b000111011011: colour_data = 24'b111111110000000010010110;
		12'b000111011100: colour_data = 24'b111111110000000010010110;
		12'b000111011101: colour_data = 24'b001000100010001011001100;
		12'b000111011110: colour_data = 24'b001000100010001011001100;
		12'b000111011111: colour_data = 24'b111111110000000010010110;
		12'b000111100000: colour_data = 24'b111111110000000010010110;
		12'b000111100001: colour_data = 24'b111111110000000010010110;
		12'b000111100010: colour_data = 24'b111111110000000010010110;
		12'b000111100011: colour_data = 24'b111111110000000010010110;
		12'b000111100100: colour_data = 24'b111111110000000010010110;

		12'b001000000000: colour_data = 24'b111111110000000010010110;
		12'b001000000001: colour_data = 24'b111111110000000010010110;
		12'b001000000010: colour_data = 24'b111111110000000010010110;
		12'b001000000011: colour_data = 24'b111111110000000010010110;
		12'b001000000100: colour_data = 24'b111111110000000010010110;
		12'b001000000101: colour_data = 24'b111111110000000010010110;
		12'b001000000110: colour_data = 24'b111111110000000010010110;
		12'b001000000111: colour_data = 24'b111111110000000010010110;
		12'b001000001000: colour_data = 24'b111111110000000010010110;
		12'b001000001001: colour_data = 24'b111111110000000010010110;
		12'b001000001010: colour_data = 24'b111111110000000010010110;
		12'b001000001011: colour_data = 24'b111111110000000010010110;
		12'b001000001100: colour_data = 24'b111111110000000010010110;
		12'b001000001101: colour_data = 24'b111111110000000010010110;
		12'b001000001110: colour_data = 24'b001000100010001011001100;
		12'b001000001111: colour_data = 24'b001000100010001011001100;
		12'b001000010000: colour_data = 24'b001000100010001011001100;
		12'b001000010001: colour_data = 24'b001000100010001011001100;
		12'b001000010010: colour_data = 24'b101101000110110001001000;
		12'b001000010011: colour_data = 24'b111111001011010010010000;
		12'b001000010100: colour_data = 24'b010001000100010011101110;
		12'b001000010101: colour_data = 24'b010001000100010011101110;
		12'b001000010110: colour_data = 24'b010001000100010011101110;
		12'b001000010111: colour_data = 24'b010001000100010011101110;
		12'b001000011000: colour_data = 24'b010001000100010011101110;
		12'b001000011001: colour_data = 24'b011001100110011011101110;
		12'b001000011010: colour_data = 24'b100010001000100011101110;
		12'b001000011011: colour_data = 24'b001000100010001011001100;
		12'b001000011100: colour_data = 24'b001000100010001011001100;
		12'b001000011101: colour_data = 24'b001000100010001011001100;
		12'b001000011110: colour_data = 24'b001000100010001011001100;
		12'b001000011111: colour_data = 24'b111111110000000010010110;
		12'b001000100000: colour_data = 24'b111111110000000010010110;
		12'b001000100001: colour_data = 24'b111111110000000010010110;
		12'b001000100010: colour_data = 24'b111111110000000010010110;
		12'b001000100011: colour_data = 24'b111111110000000010010110;
		12'b001000100100: colour_data = 24'b111111110000000010010110;

		12'b001001000000: colour_data = 24'b111111110000000010010110;
		12'b001001000001: colour_data = 24'b111111110000000010010110;
		12'b001001000010: colour_data = 24'b111111110000000010010110;
		12'b001001000011: colour_data = 24'b111111110000000010010110;
		12'b001001000100: colour_data = 24'b111111110000000010010110;
		12'b001001000101: colour_data = 24'b111111110000000010010110;
		12'b001001000110: colour_data = 24'b111111110000000010010110;
		12'b001001000111: colour_data = 24'b111111110000000010010110;
		12'b001001001000: colour_data = 24'b111111110000000010010110;
		12'b001001001001: colour_data = 24'b111111110000000010010110;
		12'b001001001010: colour_data = 24'b111111110000000010010110;
		12'b001001001011: colour_data = 24'b111111110000000010010110;
		12'b001001001100: colour_data = 24'b111111110000000010010110;
		12'b001001001101: colour_data = 24'b111111110000000010010110;
		12'b001001001110: colour_data = 24'b111111110000000010010110;
		12'b001001001111: colour_data = 24'b001000100010001011001100;
		12'b001001010000: colour_data = 24'b001000100010001011001100;
		12'b001001010001: colour_data = 24'b001000100010001011001100;
		12'b001001010010: colour_data = 24'b111111001011010010010000;
		12'b001001010011: colour_data = 24'b111111001011010010010000;
		12'b001001010100: colour_data = 24'b101101000110110001001000;
		12'b001001010101: colour_data = 24'b010001000100010011101110;
		12'b001001010110: colour_data = 24'b010001000100010011101110;
		12'b001001010111: colour_data = 24'b010001000100010011101110;
		12'b001001011000: colour_data = 24'b010001000100010011101110;
		12'b001001011001: colour_data = 24'b010001000100010011101110;
		12'b001001011010: colour_data = 24'b011001100110011011101110;
		12'b001001011011: colour_data = 24'b100010001000100011101110;
		12'b001001011100: colour_data = 24'b001000100010001011001100;
		12'b001001011101: colour_data = 24'b001000100010001011001100;
		12'b001001011110: colour_data = 24'b001000100010001011001100;
		12'b001001011111: colour_data = 24'b111111110000000010010110;
		12'b001001100000: colour_data = 24'b111111110000000010010110;
		12'b001001100001: colour_data = 24'b111111110000000010010110;
		12'b001001100010: colour_data = 24'b111111110000000010010110;
		12'b001001100011: colour_data = 24'b111111110000000010010110;
		12'b001001100100: colour_data = 24'b111111110000000010010110;

		12'b001010000000: colour_data = 24'b111111110000000010010110;
		12'b001010000001: colour_data = 24'b111111110000000010010110;
		12'b001010000010: colour_data = 24'b111111110000000010010110;
		12'b001010000011: colour_data = 24'b111111110000000010010110;
		12'b001010000100: colour_data = 24'b111111110000000010010110;
		12'b001010000101: colour_data = 24'b111111110000000010010110;
		12'b001010000110: colour_data = 24'b111111110000000010010110;
		12'b001010000111: colour_data = 24'b111111110000000010010110;
		12'b001010001000: colour_data = 24'b111111110000000010010110;
		12'b001010001001: colour_data = 24'b111111110000000010010110;
		12'b001010001010: colour_data = 24'b111111110000000010010110;
		12'b001010001011: colour_data = 24'b111111110000000010010110;
		12'b001010001100: colour_data = 24'b111111110000000010010110;
		12'b001010001101: colour_data = 24'b111111110000000010010110;
		12'b001010001110: colour_data = 24'b111111110000000010010110;
		12'b001010001111: colour_data = 24'b001000100010001011001100;
		12'b001010010000: colour_data = 24'b001000100010001011001100;
		12'b001010010001: colour_data = 24'b001000100010001011001100;
		12'b001010010010: colour_data = 24'b111111001011010010010000;
		12'b001010010011: colour_data = 24'b111111001011010010010000;
		12'b001010010100: colour_data = 24'b111111001011010010010000;
		12'b001010010101: colour_data = 24'b101101000110110001001000;
		12'b001010010110: colour_data = 24'b010001000100010011101110;
		12'b001010010111: colour_data = 24'b010001000100010011101110;
		12'b001010011000: colour_data = 24'b010001000100010011101110;
		12'b001010011001: colour_data = 24'b010001000100010011101110;
		12'b001010011010: colour_data = 24'b010001000100010011101110;
		12'b001010011011: colour_data = 24'b011001100110011011101110;
		12'b001010011100: colour_data = 24'b100010001000100011101110;
		12'b001010011101: colour_data = 24'b001000100010001011001100;
		12'b001010011110: colour_data = 24'b111111110000000010010110;
		12'b001010011111: colour_data = 24'b111111110000000010010110;
		12'b001010100000: colour_data = 24'b111111110000000010010110;
		12'b001010100001: colour_data = 24'b111111110000000010010110;
		12'b001010100010: colour_data = 24'b111111110000000010010110;
		12'b001010100011: colour_data = 24'b111111110000000010010110;
		12'b001010100100: colour_data = 24'b111111110000000010010110;

		12'b001011000000: colour_data = 24'b111111110000000010010110;
		12'b001011000001: colour_data = 24'b111111110000000010010110;
		12'b001011000010: colour_data = 24'b111111110000000010010110;
		12'b001011000011: colour_data = 24'b111111110000000010010110;
		12'b001011000100: colour_data = 24'b111111110000000010010110;
		12'b001011000101: colour_data = 24'b111111110000000010010110;
		12'b001011000110: colour_data = 24'b111111110000000010010110;
		12'b001011000111: colour_data = 24'b111111110000000010010110;
		12'b001011001000: colour_data = 24'b111111110000000010010110;
		12'b001011001001: colour_data = 24'b111111110000000010010110;
		12'b001011001010: colour_data = 24'b111111110000000010010110;
		12'b001011001011: colour_data = 24'b111111110000000010010110;
		12'b001011001100: colour_data = 24'b111111110000000010010110;
		12'b001011001101: colour_data = 24'b111111110000000010010110;
		12'b001011001110: colour_data = 24'b010001000100010011101110;
		12'b001011001111: colour_data = 24'b001000100010001011001100;
		12'b001011010000: colour_data = 24'b010001000100010011101110;
		12'b001011010001: colour_data = 24'b010001000100010011101110;
		12'b001011010010: colour_data = 24'b001000100010001011001100;
		12'b001011010011: colour_data = 24'b111111001011010010010000;
		12'b001011010100: colour_data = 24'b111111001011010010010000;
		12'b001011010101: colour_data = 24'b010001000100010011101110;
		12'b001011010110: colour_data = 24'b010001000100010011101110;
		12'b001011010111: colour_data = 24'b010001000100010011101110;
		12'b001011011000: colour_data = 24'b010001000100010011101110;
		12'b001011011001: colour_data = 24'b010001000100010011101110;
		12'b001011011010: colour_data = 24'b010001000100010011101110;
		12'b001011011011: colour_data = 24'b010001000100010011101110;
		12'b001011011100: colour_data = 24'b011001100110011011101110;
		12'b001011011101: colour_data = 24'b100010001000100011101110;
		12'b001011011110: colour_data = 24'b111111110000000010010110;
		12'b001011011111: colour_data = 24'b111111110000000010010110;
		12'b001011100000: colour_data = 24'b111111110000000010010110;
		12'b001011100001: colour_data = 24'b111111110000000010010110;
		12'b001011100010: colour_data = 24'b111111110000000010010110;
		12'b001011100011: colour_data = 24'b111111110000000010010110;
		12'b001011100100: colour_data = 24'b111111110000000010010110;

		12'b001100000000: colour_data = 24'b111111110000000010010110;
		12'b001100000001: colour_data = 24'b111111110000000010010110;
		12'b001100000010: colour_data = 24'b111111110000000010010110;
		12'b001100000011: colour_data = 24'b111111110000000010010110;
		12'b001100000100: colour_data = 24'b111111110000000010010110;
		12'b001100000101: colour_data = 24'b111111110000000010010110;
		12'b001100000110: colour_data = 24'b111111110000000010010110;
		12'b001100000111: colour_data = 24'b111111110000000010010110;
		12'b001100001000: colour_data = 24'b111111110000000010010110;
		12'b001100001001: colour_data = 24'b111111110000000010010110;
		12'b001100001010: colour_data = 24'b111111110000000010010110;
		12'b001100001011: colour_data = 24'b111111110000000010010110;
		12'b001100001100: colour_data = 24'b010001000100010011101110;
		12'b001100001101: colour_data = 24'b010001000100010011101110;
		12'b001100001110: colour_data = 24'b001000100010001011001100;
		12'b001100001111: colour_data = 24'b010001000100010011101110;
		12'b001100010000: colour_data = 24'b010001000100010011101110;
		12'b001100010001: colour_data = 24'b010001000100010011101110;
		12'b001100010010: colour_data = 24'b010001000100010011101110;
		12'b001100010011: colour_data = 24'b111111001011010010010000;
		12'b001100010100: colour_data = 24'b010001000100010011101110;
		12'b001100010101: colour_data = 24'b010001000100010011101110;
		12'b001100010110: colour_data = 24'b010001000100010011101110;
		12'b001100010111: colour_data = 24'b010001000100010011101110;
		12'b001100011000: colour_data = 24'b010001000100010011101110;
		12'b001100011001: colour_data = 24'b010001000100010011101110;
		12'b001100011010: colour_data = 24'b010001000100010011101110;
		12'b001100011011: colour_data = 24'b010001000100010011101110;
		12'b001100011100: colour_data = 24'b010001000100010011101110;
		12'b001100011101: colour_data = 24'b100010001000100011101110;
		12'b001100011110: colour_data = 24'b111111110000000010010110;
		12'b001100011111: colour_data = 24'b111111110000000010010110;
		12'b001100100000: colour_data = 24'b111111110000000010010110;
		12'b001100100001: colour_data = 24'b111111110000000010010110;
		12'b001100100010: colour_data = 24'b111111110000000010010110;
		12'b001100100011: colour_data = 24'b111111110000000010010110;
		12'b001100100100: colour_data = 24'b111111110000000010010110;

		12'b001101000000: colour_data = 24'b111111110000000010010110;
		12'b001101000001: colour_data = 24'b111111110000000010010110;
		12'b001101000010: colour_data = 24'b111111110000000010010110;
		12'b001101000011: colour_data = 24'b111111110000000010010110;
		12'b001101000100: colour_data = 24'b111111110000000010010110;
		12'b001101000101: colour_data = 24'b111111110000000010010110;
		12'b001101000110: colour_data = 24'b111111110000000010010110;
		12'b001101000111: colour_data = 24'b111111110000000010010110;
		12'b001101001000: colour_data = 24'b111111110000000010010110;
		12'b001101001001: colour_data = 24'b111111110000000010010110;
		12'b001101001010: colour_data = 24'b010001000100010011101110;
		12'b001101001011: colour_data = 24'b010001000100010011101110;
		12'b001101001100: colour_data = 24'b001000100010001011001100;
		12'b001101001101: colour_data = 24'b001000100010001011001100;
		12'b001101001110: colour_data = 24'b010001000100010011101110;
		12'b001101001111: colour_data = 24'b010001000100010011101110;
		12'b001101010000: colour_data = 24'b010001000100010011101110;
		12'b001101010001: colour_data = 24'b010001000100010011101110;
		12'b001101010010: colour_data = 24'b010001000100010011101110;
		12'b001101010011: colour_data = 24'b010001000100010011101110;
		12'b001101010100: colour_data = 24'b010001000100010011101110;
		12'b001101010101: colour_data = 24'b010001000100010011101110;
		12'b001101010110: colour_data = 24'b010001000100010011101110;
		12'b001101010111: colour_data = 24'b011001100110011011101110;
		12'b001101011000: colour_data = 24'b111111001111110011111100;
		12'b001101011001: colour_data = 24'b011001100110011011101110;
		12'b001101011010: colour_data = 24'b010001000100010011101110;
		12'b001101011011: colour_data = 24'b010001000100010011101110;
		12'b001101011100: colour_data = 24'b010001000100010011101110;
		12'b001101011101: colour_data = 24'b011001100110011011101110;
		12'b001101011110: colour_data = 24'b100010001000100011101110;
		12'b001101011111: colour_data = 24'b111111110000000010010110;
		12'b001101100000: colour_data = 24'b111111110000000010010110;
		12'b001101100001: colour_data = 24'b111111110000000010010110;
		12'b001101100010: colour_data = 24'b111111110000000010010110;
		12'b001101100011: colour_data = 24'b111111110000000010010110;
		12'b001101100100: colour_data = 24'b111111110000000010010110;

		12'b001110000000: colour_data = 24'b111111110000000010010110;
		12'b001110000001: colour_data = 24'b111111110000000010010110;
		12'b001110000010: colour_data = 24'b111111110000000010010110;
		12'b001110000011: colour_data = 24'b111111110000000010010110;
		12'b001110000100: colour_data = 24'b111111110000000010010110;
		12'b001110000101: colour_data = 24'b111111110000000010010110;
		12'b001110000110: colour_data = 24'b111111110000000010010110;
		12'b001110000111: colour_data = 24'b111111110000000010010110;
		12'b001110001000: colour_data = 24'b111111110000000010010110;
		12'b001110001001: colour_data = 24'b010001000100010011101110;
		12'b001110001010: colour_data = 24'b001000100010001011001100;
		12'b001110001011: colour_data = 24'b001000100010001011001100;
		12'b001110001100: colour_data = 24'b001000100010001011001100;
		12'b001110001101: colour_data = 24'b001000100010001011001100;
		12'b001110001110: colour_data = 24'b010001000100010011101110;
		12'b001110001111: colour_data = 24'b011001100110011011101110;
		12'b001110010000: colour_data = 24'b010001000100010011101110;
		12'b001110010001: colour_data = 24'b010001000100010011101110;
		12'b001110010010: colour_data = 24'b010001000100010011101110;
		12'b001110010011: colour_data = 24'b010001000100010011101110;
		12'b001110010100: colour_data = 24'b010001000100010011101110;
		12'b001110010101: colour_data = 24'b010001000100010011101110;
		12'b001110010110: colour_data = 24'b011001100110011011101110;
		12'b001110010111: colour_data = 24'b111111001111110011111100;
		12'b001110011000: colour_data = 24'b111111001111110011111100;
		12'b001110011001: colour_data = 24'b111111001111110011111100;
		12'b001110011010: colour_data = 24'b011001100110011011101110;
		12'b001110011011: colour_data = 24'b010001000100010011101110;
		12'b001110011100: colour_data = 24'b010001000100010011101110;
		12'b001110011101: colour_data = 24'b011001100110011011101110;
		12'b001110011110: colour_data = 24'b100010001000100011101110;
		12'b001110011111: colour_data = 24'b111111110000000010010110;
		12'b001110100000: colour_data = 24'b111111110000000010010110;
		12'b001110100001: colour_data = 24'b111111110000000010010110;
		12'b001110100010: colour_data = 24'b111111110000000010010110;
		12'b001110100011: colour_data = 24'b111111110000000010010110;
		12'b001110100100: colour_data = 24'b111111110000000010010110;

		12'b001111000000: colour_data = 24'b111111110000000010010110;
		12'b001111000001: colour_data = 24'b111111110000000010010110;
		12'b001111000010: colour_data = 24'b111111110000000010010110;
		12'b001111000011: colour_data = 24'b111111110000000010010110;
		12'b001111000100: colour_data = 24'b111111110000000010010110;
		12'b001111000101: colour_data = 24'b111111110000000010010110;
		12'b001111000110: colour_data = 24'b111111110000000010010110;
		12'b001111000111: colour_data = 24'b111111110000000010010110;
		12'b001111001000: colour_data = 24'b010001000100010011101110;
		12'b001111001001: colour_data = 24'b001000100010001011001100;
		12'b001111001010: colour_data = 24'b001000100010001011001100;
		12'b001111001011: colour_data = 24'b001000100010001011001100;
		12'b001111001100: colour_data = 24'b001000100010001011001100;
		12'b001111001101: colour_data = 24'b001000100010001011001100;
		12'b001111001110: colour_data = 24'b010001000100010011101110;
		12'b001111001111: colour_data = 24'b011001100110011011101110;
		12'b001111010000: colour_data = 24'b010001000100010011101110;
		12'b001111010001: colour_data = 24'b010001000100010011101110;
		12'b001111010010: colour_data = 24'b010001000100010011101110;
		12'b001111010011: colour_data = 24'b010001000100010011101110;
		12'b001111010100: colour_data = 24'b010001000100010011101110;
		12'b001111010101: colour_data = 24'b010001000100010011101110;
		12'b001111010110: colour_data = 24'b100010001000100011101110;
		12'b001111010111: colour_data = 24'b111111001111110011111100;
		12'b001111011000: colour_data = 24'b111111001111110011111100;
		12'b001111011001: colour_data = 24'b111111001111110011111100;
		12'b001111011010: colour_data = 24'b000000000000000000000000;
		12'b001111011011: colour_data = 24'b011001100110011011101110;
		12'b001111011100: colour_data = 24'b010001000100010011101110;
		12'b001111011101: colour_data = 24'b011001100110011011101110;
		12'b001111011110: colour_data = 24'b000000000000000000000000;
		12'b001111011111: colour_data = 24'b111111110000000010010110;
		12'b001111100000: colour_data = 24'b111111110000000010010110;
		12'b001111100001: colour_data = 24'b111111110000000010010110;
		12'b001111100010: colour_data = 24'b111111110000000010010110;
		12'b001111100011: colour_data = 24'b111111110000000010010110;
		12'b001111100100: colour_data = 24'b111111110000000010010110;

		12'b010000000000: colour_data = 24'b111111110000000010010110;
		12'b010000000001: colour_data = 24'b111111110000000010010110;
		12'b010000000010: colour_data = 24'b111111110000000010010110;
		12'b010000000011: colour_data = 24'b111111110000000010010110;
		12'b010000000100: colour_data = 24'b111111110000000010010110;
		12'b010000000101: colour_data = 24'b111111110000000010010110;
		12'b010000000110: colour_data = 24'b111111110000000010010110;
		12'b010000000111: colour_data = 24'b010001000100010011101110;
		12'b010000001000: colour_data = 24'b001000100010001011001100;
		12'b010000001001: colour_data = 24'b001000100010001011001100;
		12'b010000001010: colour_data = 24'b001000100010001011001100;
		12'b010000001011: colour_data = 24'b001000100010001011001100;
		12'b010000001100: colour_data = 24'b001000100010001011001100;
		12'b010000001101: colour_data = 24'b001000100010001011001100;
		12'b010000001110: colour_data = 24'b010001000100010011101110;
		12'b010000001111: colour_data = 24'b011001100110011011101110;
		12'b010000010000: colour_data = 24'b010001000100010011101110;
		12'b010000010001: colour_data = 24'b010001000100010011101110;
		12'b010000010010: colour_data = 24'b010001000100010011101110;
		12'b010000010011: colour_data = 24'b010001000100010011101110;
		12'b010000010100: colour_data = 24'b010001000100010011101110;
		12'b010000010101: colour_data = 24'b010001000100010011101110;
		12'b010000010110: colour_data = 24'b100010001000100011101110;
		12'b010000010111: colour_data = 24'b111111001111110011111100;
		12'b010000011000: colour_data = 24'b111111001111110011111100;
		12'b010000011001: colour_data = 24'b111111001111110011111100;
		12'b010000011010: colour_data = 24'b000000000000000000000000;
		12'b010000011011: colour_data = 24'b000000000000000000000000;
		12'b010000011100: colour_data = 24'b011001100110011011101110;
		12'b010000011101: colour_data = 24'b000000000000000000000000;
		12'b010000011110: colour_data = 24'b000000000000000000000000;
		12'b010000011111: colour_data = 24'b111111110000000010010110;
		12'b010000100000: colour_data = 24'b111111110000000010010110;
		12'b010000100001: colour_data = 24'b111111110000000010010110;
		12'b010000100010: colour_data = 24'b111111110000000010010110;
		12'b010000100011: colour_data = 24'b111111110000000010010110;
		12'b010000100100: colour_data = 24'b111111110000000010010110;

		12'b010001000000: colour_data = 24'b111111110000000010010110;
		12'b010001000001: colour_data = 24'b111111110000000010010110;
		12'b010001000010: colour_data = 24'b111111110000000010010110;
		12'b010001000011: colour_data = 24'b111111110000000010010110;
		12'b010001000100: colour_data = 24'b111111110000000010010110;
		12'b010001000101: colour_data = 24'b111111110000000010010110;
		12'b010001000110: colour_data = 24'b111111110000000010010110;
		12'b010001000111: colour_data = 24'b111111110000000010010110;
		12'b010001001000: colour_data = 24'b111111110000000010010110;
		12'b010001001001: colour_data = 24'b111111110000000010010110;
		12'b010001001010: colour_data = 24'b111111110000000010010110;
		12'b010001001011: colour_data = 24'b111111110000000010010110;
		12'b010001001100: colour_data = 24'b001000100010001011001100;
		12'b010001001101: colour_data = 24'b001000100010001011001100;
		12'b010001001110: colour_data = 24'b010001000100010011101110;
		12'b010001001111: colour_data = 24'b011001100110011011101110;
		12'b010001010000: colour_data = 24'b010001000100010011101110;
		12'b010001010001: colour_data = 24'b010001000100010011101110;
		12'b010001010010: colour_data = 24'b010001000100010011101110;
		12'b010001010011: colour_data = 24'b010001000100010011101110;
		12'b010001010100: colour_data = 24'b010001000100010011101110;
		12'b010001010101: colour_data = 24'b010001000100010011101110;
		12'b010001010110: colour_data = 24'b100010001000100011101110;
		12'b010001010111: colour_data = 24'b111111001111110011111100;
		12'b010001011000: colour_data = 24'b111111001111110011111100;
		12'b010001011001: colour_data = 24'b111111001111110011111100;
		12'b010001011010: colour_data = 24'b000000000000000000000000;
		12'b010001011011: colour_data = 24'b000000000000000000000000;
		12'b010001011100: colour_data = 24'b011001100110011011101110;
		12'b010001011101: colour_data = 24'b000000000000000000000000;
		12'b010001011110: colour_data = 24'b000000000000000000000000;
		12'b010001011111: colour_data = 24'b111111110000000010010110;
		12'b010001100000: colour_data = 24'b111111110000000010010110;
		12'b010001100001: colour_data = 24'b111111110000000010010110;
		12'b010001100010: colour_data = 24'b111111110000000010010110;
		12'b010001100011: colour_data = 24'b111111110000000010010110;
		12'b010001100100: colour_data = 24'b111111110000000010010110;

		12'b010010000000: colour_data = 24'b111111110000000010010110;
		12'b010010000001: colour_data = 24'b111111110000000010010110;
		12'b010010000010: colour_data = 24'b111111110000000010010110;
		12'b010010000011: colour_data = 24'b111111110000000010010110;
		12'b010010000100: colour_data = 24'b111111110000000010010110;
		12'b010010000101: colour_data = 24'b111111110000000010010110;
		12'b010010000110: colour_data = 24'b111111110000000010010110;
		12'b010010000111: colour_data = 24'b111111110000000010010110;
		12'b010010001000: colour_data = 24'b111111110000000010010110;
		12'b010010001001: colour_data = 24'b111111110000000010010110;
		12'b010010001010: colour_data = 24'b111111110000000010010110;
		12'b010010001011: colour_data = 24'b111111110000000010010110;
		12'b010010001100: colour_data = 24'b111111110000000010010110;
		12'b010010001101: colour_data = 24'b111111110000000010010110;
		12'b010010001110: colour_data = 24'b001000100010001011001100;
		12'b010010001111: colour_data = 24'b010001000100010011101110;
		12'b010010010000: colour_data = 24'b011001100110011011101110;
		12'b010010010001: colour_data = 24'b010001000100010011101110;
		12'b010010010010: colour_data = 24'b010001000100010011101110;
		12'b010010010011: colour_data = 24'b010001000100010011101110;
		12'b010010010100: colour_data = 24'b010001000100010011101110;
		12'b010010010101: colour_data = 24'b010001000100010011101110;
		12'b010010010110: colour_data = 24'b011001100110011011101110;
		12'b010010010111: colour_data = 24'b111111001111110011111100;
		12'b010010011000: colour_data = 24'b111111001111110011111100;
		12'b010010011001: colour_data = 24'b111111001111110011111100;
		12'b010010011010: colour_data = 24'b000000000000000000000000;
		12'b010010011011: colour_data = 24'b000000000000000000000000;
		12'b010010011100: colour_data = 24'b111111001111110011111100;
		12'b010010011101: colour_data = 24'b101101001011010010110100;
		12'b010010011110: colour_data = 24'b000000000000000000000000;
		12'b010010011111: colour_data = 24'b111111110000000010010110;
		12'b010010100000: colour_data = 24'b111111110000000010010110;
		12'b010010100001: colour_data = 24'b111111110000000010010110;
		12'b010010100010: colour_data = 24'b111111110000000010010110;
		12'b010010100011: colour_data = 24'b111111110000000010010110;
		12'b010010100100: colour_data = 24'b111111110000000010010110;

		12'b010011000000: colour_data = 24'b111111110000000010010110;
		12'b010011000001: colour_data = 24'b111111110000000010010110;
		12'b010011000010: colour_data = 24'b111111110000000010010110;
		12'b010011000011: colour_data = 24'b111111110000000010010110;
		12'b010011000100: colour_data = 24'b111111110000000010010110;
		12'b010011000101: colour_data = 24'b111111110000000010010110;
		12'b010011000110: colour_data = 24'b111111110000000010010110;
		12'b010011000111: colour_data = 24'b111111110000000010010110;
		12'b010011001000: colour_data = 24'b111111110000000010010110;
		12'b010011001001: colour_data = 24'b111111110000000010010110;
		12'b010011001010: colour_data = 24'b111111110000000010010110;
		12'b010011001011: colour_data = 24'b111111110000000010010110;
		12'b010011001100: colour_data = 24'b010001000100010011101110;
		12'b010011001101: colour_data = 24'b010001000100010011101110;
		12'b010011001110: colour_data = 24'b001000100010001011001100;
		12'b010011001111: colour_data = 24'b010001000100010011101110;
		12'b010011010000: colour_data = 24'b011001100110011011101110;
		12'b010011010001: colour_data = 24'b010001000100010011101110;
		12'b010011010010: colour_data = 24'b010001000100010011101110;
		12'b010011010011: colour_data = 24'b010001000100010011101110;
		12'b010011010100: colour_data = 24'b101101000110110001001000;
		12'b010011010101: colour_data = 24'b101101000110110001001000;
		12'b010011010110: colour_data = 24'b101101000110110001001000;
		12'b010011010111: colour_data = 24'b011001100110011011101110;
		12'b010011011000: colour_data = 24'b111111001111110011111100;
		12'b010011011001: colour_data = 24'b111111001111110011111100;
		12'b010011011010: colour_data = 24'b111111001111110011111100;
		12'b010011011011: colour_data = 24'b111111001111110011111100;
		12'b010011011100: colour_data = 24'b101101001011010010110100;
		12'b010011011101: colour_data = 24'b000000000000000000000000;
		12'b010011011110: colour_data = 24'b101101001011010010110100;
		12'b010011011111: colour_data = 24'b111111110000000010010110;
		12'b010011100000: colour_data = 24'b111111110000000010010110;
		12'b010011100001: colour_data = 24'b111111110000000010010110;
		12'b010011100010: colour_data = 24'b111111110000000010010110;
		12'b010011100011: colour_data = 24'b111111110000000010010110;
		12'b010011100100: colour_data = 24'b111111110000000010010110;

		12'b010100000000: colour_data = 24'b111111110000000010010110;
		12'b010100000001: colour_data = 24'b111111110000000010010110;
		12'b010100000010: colour_data = 24'b111111110000000010010110;
		12'b010100000011: colour_data = 24'b111111110000000010010110;
		12'b010100000100: colour_data = 24'b111111110000000010010110;
		12'b010100000101: colour_data = 24'b111111110000000010010110;
		12'b010100000110: colour_data = 24'b111111110000000010010110;
		12'b010100000111: colour_data = 24'b111111110000000010010110;
		12'b010100001000: colour_data = 24'b111111110000000010010110;
		12'b010100001001: colour_data = 24'b111111110000000010010110;
		12'b010100001010: colour_data = 24'b010001000100010011101110;
		12'b010100001011: colour_data = 24'b010001000100010011101110;
		12'b010100001100: colour_data = 24'b001000100010001011001100;
		12'b010100001101: colour_data = 24'b001000100010001011001100;
		12'b010100001110: colour_data = 24'b001000100010001011001100;
		12'b010100001111: colour_data = 24'b001000100010001011001100;
		12'b010100010000: colour_data = 24'b010001000100010011101110;
		12'b010100010001: colour_data = 24'b011001100110011011101110;
		12'b010100010010: colour_data = 24'b010001000100010011101110;
		12'b010100010011: colour_data = 24'b101101000110110001001000;
		12'b010100010100: colour_data = 24'b111111001011010010010000;
		12'b010100010101: colour_data = 24'b111111001011010010010000;
		12'b010100010110: colour_data = 24'b111111001011010010010000;
		12'b010100010111: colour_data = 24'b101101000110110001001000;
		12'b010100011000: colour_data = 24'b011001100110011011101110;
		12'b010100011001: colour_data = 24'b111111001111110011111100;
		12'b010100011010: colour_data = 24'b111111001111110011111100;
		12'b010100011011: colour_data = 24'b111111001011010010010000;
		12'b010100011100: colour_data = 24'b000000000000000000000000;
		12'b010100011101: colour_data = 24'b000000000000000000000000;
		12'b010100011110: colour_data = 24'b000000000000000000000000;
		12'b010100011111: colour_data = 24'b111111110000000010010110;
		12'b010100100000: colour_data = 24'b111111110000000010010110;
		12'b010100100001: colour_data = 24'b111111110000000010010110;
		12'b010100100010: colour_data = 24'b111111110000000010010110;
		12'b010100100011: colour_data = 24'b111111110000000010010110;
		12'b010100100100: colour_data = 24'b111111110000000010010110;

		12'b010101000000: colour_data = 24'b111111110000000010010110;
		12'b010101000001: colour_data = 24'b111111110000000010010110;
		12'b010101000010: colour_data = 24'b111111110000000010010110;
		12'b010101000011: colour_data = 24'b111111110000000010010110;
		12'b010101000100: colour_data = 24'b111111110000000010010110;
		12'b010101000101: colour_data = 24'b111111110000000010010110;
		12'b010101000110: colour_data = 24'b111111110000000010010110;
		12'b010101000111: colour_data = 24'b111111110000000010010110;
		12'b010101001000: colour_data = 24'b111111110000000010010110;
		12'b010101001001: colour_data = 24'b010001000100010011101110;
		12'b010101001010: colour_data = 24'b001000100010001011001100;
		12'b010101001011: colour_data = 24'b001000100010001011001100;
		12'b010101001100: colour_data = 24'b001000100010001011001100;
		12'b010101001101: colour_data = 24'b001000100010001011001100;
		12'b010101001110: colour_data = 24'b001000100010001011001100;
		12'b010101001111: colour_data = 24'b001000100010001011001100;
		12'b010101010000: colour_data = 24'b001000100010001011001100;
		12'b010101010001: colour_data = 24'b010001000100010011101110;
		12'b010101010010: colour_data = 24'b011001100110011011101110;
		12'b010101010011: colour_data = 24'b101101000110110001001000;
		12'b010101010100: colour_data = 24'b111111001011010010010000;
		12'b010101010101: colour_data = 24'b111111001011010010010000;
		12'b010101010110: colour_data = 24'b111111001011010010010000;
		12'b010101010111: colour_data = 24'b111111001011010010010000;
		12'b010101011000: colour_data = 24'b111111001011010010010000;
		12'b010101011001: colour_data = 24'b111111001011010010010000;
		12'b010101011010: colour_data = 24'b111111001011010010010000;
		12'b010101011011: colour_data = 24'b111111001011010010010000;
		12'b010101011100: colour_data = 24'b111111001011010010010000;
		12'b010101011101: colour_data = 24'b100100001001000010010000;
		12'b010101011110: colour_data = 24'b100100001001000010010000;
		12'b010101011111: colour_data = 24'b111111110000000010010110;
		12'b010101100000: colour_data = 24'b111111110000000010010110;
		12'b010101100001: colour_data = 24'b111111110000000010010110;
		12'b010101100010: colour_data = 24'b111111110000000010010110;
		12'b010101100011: colour_data = 24'b111111110000000010010110;
		12'b010101100100: colour_data = 24'b111111110000000010010110;

		12'b010110000000: colour_data = 24'b111111110000000010010110;
		12'b010110000001: colour_data = 24'b111111110000000010010110;
		12'b010110000010: colour_data = 24'b111111110000000010010110;
		12'b010110000011: colour_data = 24'b111111110000000010010110;
		12'b010110000100: colour_data = 24'b111111110000000010010110;
		12'b010110000101: colour_data = 24'b111111110000000010010110;
		12'b010110000110: colour_data = 24'b111111110000000010010110;
		12'b010110000111: colour_data = 24'b111111110000000010010110;
		12'b010110001000: colour_data = 24'b111111110000000010010110;
		12'b010110001001: colour_data = 24'b010001000100010011101110;
		12'b010110001010: colour_data = 24'b001000100010001011001100;
		12'b010110001011: colour_data = 24'b001000100010001011001100;
		12'b010110001100: colour_data = 24'b001000100010001011001100;
		12'b010110001101: colour_data = 24'b001000100010001011001100;
		12'b010110001110: colour_data = 24'b001000100010001011001100;
		12'b010110001111: colour_data = 24'b001000100010001011001100;
		12'b010110010000: colour_data = 24'b001000100010001011001100;
		12'b010110010001: colour_data = 24'b001000100010001011001100;
		12'b010110010010: colour_data = 24'b010001000100010011101110;
		12'b010110010011: colour_data = 24'b010001000100010011101110;
		12'b010110010100: colour_data = 24'b101101000110110001001000;
		12'b010110010101: colour_data = 24'b111111001011010010010000;
		12'b010110010110: colour_data = 24'b111111001011010010010000;
		12'b010110010111: colour_data = 24'b111111001011010010010000;
		12'b010110011000: colour_data = 24'b111111001011010010010000;
		12'b010110011001: colour_data = 24'b111111001011010010010000;
		12'b010110011010: colour_data = 24'b101101000110110001001000;
		12'b010110011011: colour_data = 24'b101101000110110001001000;
		12'b010110011100: colour_data = 24'b101101001011010010110100;
		12'b010110011101: colour_data = 24'b100100001001000010010000;
		12'b010110011110: colour_data = 24'b100100001001000010010000;
		12'b010110011111: colour_data = 24'b101101001011010010110100;
		12'b010110100000: colour_data = 24'b111111110000000010010110;
		12'b010110100001: colour_data = 24'b111111110000000010010110;
		12'b010110100010: colour_data = 24'b111111110000000010010110;
		12'b010110100011: colour_data = 24'b111111110000000010010110;
		12'b010110100100: colour_data = 24'b111111110000000010010110;

		12'b010111000000: colour_data = 24'b111111110000000010010110;
		12'b010111000001: colour_data = 24'b111111110000000010010110;
		12'b010111000010: colour_data = 24'b111111110000000010010110;
		12'b010111000011: colour_data = 24'b111111110000000010010110;
		12'b010111000100: colour_data = 24'b111111110000000010010110;
		12'b010111000101: colour_data = 24'b111111110000000010010110;
		12'b010111000110: colour_data = 24'b111111110000000010010110;
		12'b010111000111: colour_data = 24'b111111110000000010010110;
		12'b010111001000: colour_data = 24'b010001000100010011101110;
		12'b010111001001: colour_data = 24'b001000100010001011001100;
		12'b010111001010: colour_data = 24'b001000100010001011001100;
		12'b010111001011: colour_data = 24'b111111001011010010010000;
		12'b010111001100: colour_data = 24'b111111001011010010010000;
		12'b010111001101: colour_data = 24'b111111001011010010010000;
		12'b010111001110: colour_data = 24'b111111001011010010010000;
		12'b010111001111: colour_data = 24'b111111001011010010010000;
		12'b010111010000: colour_data = 24'b111111001011010010010000;
		12'b010111010001: colour_data = 24'b001000100010001011001100;
		12'b010111010010: colour_data = 24'b001000100010001011001100;
		12'b010111010011: colour_data = 24'b001000100010001011001100;
		12'b010111010100: colour_data = 24'b010001000100010011101110;
		12'b010111010101: colour_data = 24'b101101000110110001001000;
		12'b010111010110: colour_data = 24'b101101000110110001001000;
		12'b010111010111: colour_data = 24'b101101000110110001001000;
		12'b010111011000: colour_data = 24'b101101000110110001001000;
		12'b010111011001: colour_data = 24'b101101000110110001001000;
		12'b010111011010: colour_data = 24'b111111110000000010010110;
		12'b010111011011: colour_data = 24'b101101001011010010110100;
		12'b010111011100: colour_data = 24'b100100001001000010010000;
		12'b010111011101: colour_data = 24'b101101001011010010110100;
		12'b010111011110: colour_data = 24'b100100001001000010010000;
		12'b010111011111: colour_data = 24'b101101001011010010110100;
		12'b010111100000: colour_data = 24'b111111110000000010010110;
		12'b010111100001: colour_data = 24'b111111110000000010010110;
		12'b010111100010: colour_data = 24'b111111110000000010010110;
		12'b010111100011: colour_data = 24'b111111110000000010010110;
		12'b010111100100: colour_data = 24'b111111110000000010010110;

		12'b011000000000: colour_data = 24'b111111110000000010010110;
		12'b011000000001: colour_data = 24'b111111110000000010010110;
		12'b011000000010: colour_data = 24'b100100001001000010010000;
		12'b011000000011: colour_data = 24'b111111001111110011111100;
		12'b011000000100: colour_data = 24'b111111001111110011111100;
		12'b011000000101: colour_data = 24'b111111001111110011111100;
		12'b011000000110: colour_data = 24'b111111001111110011111100;
		12'b011000000111: colour_data = 24'b101101001011010010110100;
		12'b011000001000: colour_data = 24'b111111001111110011111100;
		12'b011000001001: colour_data = 24'b111111001011010010010000;
		12'b011000001010: colour_data = 24'b111111001011010010010000;
		12'b011000001011: colour_data = 24'b101101000110110001001000;
		12'b011000001100: colour_data = 24'b101101000110110001001000;
		12'b011000001101: colour_data = 24'b101101000110110001001000;
		12'b011000001110: colour_data = 24'b101101000110110001001000;
		12'b011000001111: colour_data = 24'b101101000110110001001000;
		12'b011000010000: colour_data = 24'b101101000110110001001000;
		12'b011000010001: colour_data = 24'b010001000100010011101110;
		12'b011000010010: colour_data = 24'b101101000110110001001000;
		12'b011000010011: colour_data = 24'b101101000110110001001000;
		12'b011000010100: colour_data = 24'b101101000110110001001000;
		12'b011000010101: colour_data = 24'b101101000110110001001000;
		12'b011000010110: colour_data = 24'b111111001011010010010000;
		12'b011000010111: colour_data = 24'b111111110000000010010110;
		12'b011000011000: colour_data = 24'b111111110000000010010110;
		12'b011000011001: colour_data = 24'b111111110000000010010110;
		12'b011000011010: colour_data = 24'b100100001001000010010000;
		12'b011000011011: colour_data = 24'b101101001011010010110100;
		12'b011000011100: colour_data = 24'b100100001001000010010000;
		12'b011000011101: colour_data = 24'b101101001011010010110100;
		12'b011000011110: colour_data = 24'b101101001011010010110100;
		12'b011000011111: colour_data = 24'b101101001011010010110100;
		12'b011000100000: colour_data = 24'b111111110000000010010110;
		12'b011000100001: colour_data = 24'b111111110000000010010110;
		12'b011000100010: colour_data = 24'b111111110000000010010110;
		12'b011000100011: colour_data = 24'b111111110000000010010110;
		12'b011000100100: colour_data = 24'b111111110000000010010110;

		12'b011001000000: colour_data = 24'b111111110000000010010110;
		12'b011001000001: colour_data = 24'b101101001011010010110100;
		12'b011001000010: colour_data = 24'b111111001111110011111100;
		12'b011001000011: colour_data = 24'b111111001111110011111100;
		12'b011001000100: colour_data = 24'b111111001111110011111100;
		12'b011001000101: colour_data = 24'b111111001111110011111100;
		12'b011001000110: colour_data = 24'b111111001111110011111100;
		12'b011001000111: colour_data = 24'b111111001111110011111100;
		12'b011001001000: colour_data = 24'b111111001111110011111100;
		12'b011001001001: colour_data = 24'b101101000110110001001000;
		12'b011001001010: colour_data = 24'b101101000110110001001000;
		12'b011001001011: colour_data = 24'b111111110000000010010110;
		12'b011001001100: colour_data = 24'b111111110000000010010110;
		12'b011001001101: colour_data = 24'b111111110000000010010110;
		12'b011001001110: colour_data = 24'b010001000100010011101110;
		12'b011001001111: colour_data = 24'b001000100010001011001100;
		12'b011001010000: colour_data = 24'b010001000100010011101110;
		12'b011001010001: colour_data = 24'b101101000110110001001000;
		12'b011001010010: colour_data = 24'b101101000110110001001000;
		12'b011001010011: colour_data = 24'b111111001011010010010000;
		12'b011001010100: colour_data = 24'b111111001011010010010000;
		12'b011001010101: colour_data = 24'b111111001011010010010000;
		12'b011001010110: colour_data = 24'b101101000110110001001000;
		12'b011001010111: colour_data = 24'b111111001011010010010000;
		12'b011001011000: colour_data = 24'b111111001011010010010000;
		12'b011001011001: colour_data = 24'b111111001011010010010000;
		12'b011001011010: colour_data = 24'b100100001001000010010000;
		12'b011001011011: colour_data = 24'b100100001001000010010000;
		12'b011001011100: colour_data = 24'b100100001001000010010000;
		12'b011001011101: colour_data = 24'b100100001001000010010000;
		12'b011001011110: colour_data = 24'b101101001011010010110100;
		12'b011001011111: colour_data = 24'b100100001001000010010000;
		12'b011001100000: colour_data = 24'b111111110000000010010110;
		12'b011001100001: colour_data = 24'b111111110000000010010110;
		12'b011001100010: colour_data = 24'b111111110000000010010110;
		12'b011001100011: colour_data = 24'b111111110000000010010110;
		12'b011001100100: colour_data = 24'b111111110000000010010110;

		12'b011010000000: colour_data = 24'b111111110000000010010110;
		12'b011010000001: colour_data = 24'b111111001111110011111100;
		12'b011010000010: colour_data = 24'b111111001111110011111100;
		12'b011010000011: colour_data = 24'b111111001111110011111100;
		12'b011010000100: colour_data = 24'b111111001111110011111100;
		12'b011010000101: colour_data = 24'b111111001111110011111100;
		12'b011010000110: colour_data = 24'b111111001111110011111100;
		12'b011010000111: colour_data = 24'b100100001001000010010000;
		12'b011010001000: colour_data = 24'b101101001011010010110100;
		12'b011010001001: colour_data = 24'b111111110000000010010110;
		12'b011010001010: colour_data = 24'b111111110000000010010110;
		12'b011010001011: colour_data = 24'b111111110000000010010110;
		12'b011010001100: colour_data = 24'b111111110000000010010110;
		12'b011010001101: colour_data = 24'b010001000100010011101110;
		12'b011010001110: colour_data = 24'b001000100010001011001100;
		12'b011010001111: colour_data = 24'b001000100010001011001100;
		12'b011010010000: colour_data = 24'b010001000100010011101110;
		12'b011010010001: colour_data = 24'b101101000110110001001000;
		12'b011010010010: colour_data = 24'b111111001011010010010000;
		12'b011010010011: colour_data = 24'b111111001011010010010000;
		12'b011010010100: colour_data = 24'b111111001011010010010000;
		12'b011010010101: colour_data = 24'b111111001011010010010000;
		12'b011010010110: colour_data = 24'b111111001011010010010000;
		12'b011010010111: colour_data = 24'b101101000110110001001000;
		12'b011010011000: colour_data = 24'b101101000110110001001000;
		12'b011010011001: colour_data = 24'b101101000110110001001000;
		12'b011010011010: colour_data = 24'b111111110000000010010110;
		12'b011010011011: colour_data = 24'b100100001001000010010000;
		12'b011010011100: colour_data = 24'b100100001001000010010000;
		12'b011010011101: colour_data = 24'b101101001011010010110100;
		12'b011010011110: colour_data = 24'b100100001001000010010000;
		12'b011010011111: colour_data = 24'b111111110000000010010110;
		12'b011010100000: colour_data = 24'b111111110000000010010110;
		12'b011010100001: colour_data = 24'b111111110000000010010110;
		12'b011010100010: colour_data = 24'b111111110000000010010110;
		12'b011010100011: colour_data = 24'b111111110000000010010110;
		12'b011010100100: colour_data = 24'b111111110000000010010110;

		12'b011011000000: colour_data = 24'b111111110000000010010110;
		12'b011011000001: colour_data = 24'b101101001011010010110100;
		12'b011011000010: colour_data = 24'b111111001111110011111100;
		12'b011011000011: colour_data = 24'b111111001111110011111100;
		12'b011011000100: colour_data = 24'b111111001111110011111100;
		12'b011011000101: colour_data = 24'b111111001111110011111100;
		12'b011011000110: colour_data = 24'b111111001111110011111100;
		12'b011011000111: colour_data = 24'b101101001011010010110100;
		12'b011011001000: colour_data = 24'b111111110000000010010110;
		12'b011011001001: colour_data = 24'b111111110000000010010110;
		12'b011011001010: colour_data = 24'b111111110000000010010110;
		12'b011011001011: colour_data = 24'b111111110000000010010110;
		12'b011011001100: colour_data = 24'b010001000100010011101110;
		12'b011011001101: colour_data = 24'b001000100010001011001100;
		12'b011011001110: colour_data = 24'b001000100010001011001100;
		12'b011011001111: colour_data = 24'b001000100010001011001100;
		12'b011011010000: colour_data = 24'b010001000100010011101110;
		12'b011011010001: colour_data = 24'b101101000110110001001000;
		12'b011011010010: colour_data = 24'b111111001011010010010000;
		12'b011011010011: colour_data = 24'b111111001011010010010000;
		12'b011011010100: colour_data = 24'b111111001011010010010000;
		12'b011011010101: colour_data = 24'b111111001011010010010000;
		12'b011011010110: colour_data = 24'b111111001011010010010000;
		12'b011011010111: colour_data = 24'b111111110000000010010110;
		12'b011011011000: colour_data = 24'b111111110000000010010110;
		12'b011011011001: colour_data = 24'b111111110000000010010110;
		12'b011011011010: colour_data = 24'b111111110000000010010110;
		12'b011011011011: colour_data = 24'b111111110000000010010110;
		12'b011011011100: colour_data = 24'b111111110000000010010110;
		12'b011011011101: colour_data = 24'b111111110000000010010110;
		12'b011011011110: colour_data = 24'b111111110000000010010110;
		12'b011011011111: colour_data = 24'b111111110000000010010110;
		12'b011011100000: colour_data = 24'b111111110000000010010110;
		12'b011011100001: colour_data = 24'b111111110000000010010110;
		12'b011011100010: colour_data = 24'b111111110000000010010110;
		12'b011011100011: colour_data = 24'b111111110000000010010110;
		12'b011011100100: colour_data = 24'b111111110000000010010110;

		12'b011100000000: colour_data = 24'b111111110000000010010110;
		12'b011100000001: colour_data = 24'b101101001011010010110100;
		12'b011100000010: colour_data = 24'b111111001111110011111100;
		12'b011100000011: colour_data = 24'b111111001111110011111100;
		12'b011100000100: colour_data = 24'b100100001001000010010000;
		12'b011100000101: colour_data = 24'b111111001111110011111100;
		12'b011100000110: colour_data = 24'b101101001011010010110100;
		12'b011100000111: colour_data = 24'b111111110000000010010110;
		12'b011100001000: colour_data = 24'b111111110000000010010110;
		12'b011100001001: colour_data = 24'b111111110000000010010110;
		12'b011100001010: colour_data = 24'b111111110000000010010110;
		12'b011100001011: colour_data = 24'b111111110000000010010110;
		12'b011100001100: colour_data = 24'b010001000100010011101110;
		12'b011100001101: colour_data = 24'b001000100010001011001100;
		12'b011100001110: colour_data = 24'b001000100010001011001100;
		12'b011100001111: colour_data = 24'b001000100010001011001100;
		12'b011100010000: colour_data = 24'b001000100010001011001100;
		12'b011100010001: colour_data = 24'b010001000100010011101110;
		12'b011100010010: colour_data = 24'b011001100110011011101110;
		12'b011100010011: colour_data = 24'b101101000110110001001000;
		12'b011100010100: colour_data = 24'b101101000110110001001000;
		12'b011100010101: colour_data = 24'b111111001011010010010000;
		12'b011100010110: colour_data = 24'b101101000110110001001000;
		12'b011100010111: colour_data = 24'b111111110000000010010110;
		12'b011100011000: colour_data = 24'b111111110000000010010110;
		12'b011100011001: colour_data = 24'b111111110000000010010110;
		12'b011100011010: colour_data = 24'b111111110000000010010110;
		12'b011100011011: colour_data = 24'b111111110000000010010110;
		12'b011100011100: colour_data = 24'b111111110000000010010110;
		12'b011100011101: colour_data = 24'b111111110000000010010110;
		12'b011100011110: colour_data = 24'b111111110000000010010110;
		12'b011100011111: colour_data = 24'b111111110000000010010110;
		12'b011100100000: colour_data = 24'b111111110000000010010110;
		12'b011100100001: colour_data = 24'b111111110000000010010110;
		12'b011100100010: colour_data = 24'b111111000000000000000000;
		12'b011100100011: colour_data = 24'b111111000000000000000000;
		12'b011100100100: colour_data = 24'b000000000000000000000000;

		12'b011101000000: colour_data = 24'b111111110000000010010110;
		12'b011101000001: colour_data = 24'b111111110000000010010110;
		12'b011101000010: colour_data = 24'b111111001111110011111100;
		12'b011101000011: colour_data = 24'b100100001001000010010000;
		12'b011101000100: colour_data = 24'b111111001111110011111100;
		12'b011101000101: colour_data = 24'b101101001011010010110100;
		12'b011101000110: colour_data = 24'b111111110000000010010110;
		12'b011101000111: colour_data = 24'b111111110000000010010110;
		12'b011101001000: colour_data = 24'b111111110000000010010110;
		12'b011101001001: colour_data = 24'b000000000000000000000000;
		12'b011101001010: colour_data = 24'b100100000000000000000000;
		12'b011101001011: colour_data = 24'b010001000100010011101110;
		12'b011101001100: colour_data = 24'b001000100010001011001100;
		12'b011101001101: colour_data = 24'b001000100010001011001100;
		12'b011101001110: colour_data = 24'b001000100010001011001100;
		12'b011101001111: colour_data = 24'b111111110000000010010110;
		12'b011101010000: colour_data = 24'b001000100010001011001100;
		12'b011101010001: colour_data = 24'b001000100010001011001100;
		12'b011101010010: colour_data = 24'b010001000100010011101110;
		12'b011101010011: colour_data = 24'b011001100110011011101110;
		12'b011101010100: colour_data = 24'b011001100110011011101110;
		12'b011101010101: colour_data = 24'b011001100110011011101110;
		12'b011101010110: colour_data = 24'b011001100110011011101110;
		12'b011101010111: colour_data = 24'b111111110000000010010110;
		12'b011101011000: colour_data = 24'b111111110000000010010110;
		12'b011101011001: colour_data = 24'b111111110000000010010110;
		12'b011101011010: colour_data = 24'b111111110000000010010110;
		12'b011101011011: colour_data = 24'b111111110000000010010110;
		12'b011101011100: colour_data = 24'b111111110000000010010110;
		12'b011101011101: colour_data = 24'b111111110000000010010110;
		12'b011101011110: colour_data = 24'b111111110000000010010110;
		12'b011101011111: colour_data = 24'b111111110000000010010110;
		12'b011101100000: colour_data = 24'b111111110000000010010110;
		12'b011101100001: colour_data = 24'b111111000000000000000000;
		12'b011101100010: colour_data = 24'b111111000000000000000000;
		12'b011101100011: colour_data = 24'b111111000000000000000000;
		12'b011101100100: colour_data = 24'b000000000000000000000000;

		12'b011110000000: colour_data = 24'b111111110000000010010110;
		12'b011110000001: colour_data = 24'b111111110000000010010110;
		12'b011110000010: colour_data = 24'b111111110000000010010110;
		12'b011110000011: colour_data = 24'b111111110000000010010110;
		12'b011110000100: colour_data = 24'b111111110000000010010110;
		12'b011110000101: colour_data = 24'b111111110000000010010110;
		12'b011110000110: colour_data = 24'b111111110000000010010110;
		12'b011110000111: colour_data = 24'b111111110000000010010110;
		12'b011110001000: colour_data = 24'b000000000000000000000000;
		12'b011110001001: colour_data = 24'b100100000000000000000000;
		12'b011110001010: colour_data = 24'b000000000000000000000000;
		12'b011110001011: colour_data = 24'b010001000100010011101110;
		12'b011110001100: colour_data = 24'b100100000000000000000000;
		12'b011110001101: colour_data = 24'b101101001011010010110100;
		12'b011110001110: colour_data = 24'b101101001011010010110100;
		12'b011110001111: colour_data = 24'b111111110000000010010110;
		12'b011110010000: colour_data = 24'b000000000000000000000000;
		12'b011110010001: colour_data = 24'b001000100010001011001100;
		12'b011110010010: colour_data = 24'b001000100010001011001100;
		12'b011110010011: colour_data = 24'b010001000100010011101110;
		12'b011110010100: colour_data = 24'b010001000100010011101110;
		12'b011110010101: colour_data = 24'b010001000100010011101110;
		12'b011110010110: colour_data = 24'b010001000100010011101110;
		12'b011110010111: colour_data = 24'b011001100110011011101110;
		12'b011110011000: colour_data = 24'b011001100110011011101110;
		12'b011110011001: colour_data = 24'b111111110000000010010110;
		12'b011110011010: colour_data = 24'b111111110000000010010110;
		12'b011110011011: colour_data = 24'b111111110000000010010110;
		12'b011110011100: colour_data = 24'b111111110000000010010110;
		12'b011110011101: colour_data = 24'b111111110000000010010110;
		12'b011110011110: colour_data = 24'b111111110000000010010110;
		12'b011110011111: colour_data = 24'b111111000000000000000000;
		12'b011110100000: colour_data = 24'b111111000000000000000000;
		12'b011110100001: colour_data = 24'b111111000000000000000000;
		12'b011110100010: colour_data = 24'b111111000000000000000000;
		12'b011110100011: colour_data = 24'b000000000000000000000000;
		12'b011110100100: colour_data = 24'b111111110000000010010110;

		12'b011111000000: colour_data = 24'b111111110000000010010110;
		12'b011111000001: colour_data = 24'b111111110000000010010110;
		12'b011111000010: colour_data = 24'b111111110000000010010110;
		12'b011111000011: colour_data = 24'b111111110000000010010110;
		12'b011111000100: colour_data = 24'b111111110000000010010110;
		12'b011111000101: colour_data = 24'b111111110000000010010110;
		12'b011111000110: colour_data = 24'b111111110000000010010110;
		12'b011111000111: colour_data = 24'b111111110000000010010110;
		12'b011111001000: colour_data = 24'b000000000000000000000000;
		12'b011111001001: colour_data = 24'b100100000000000000000000;
		12'b011111001010: colour_data = 24'b000000000000000000000000;
		12'b011111001011: colour_data = 24'b100100000000000000000000;
		12'b011111001100: colour_data = 24'b100100000000000000000000;
		12'b011111001101: colour_data = 24'b100100000000000000000000;
		12'b011111001110: colour_data = 24'b101101001011010010110100;
		12'b011111001111: colour_data = 24'b111111110000000010010110;
		12'b011111010000: colour_data = 24'b001000100010001011001100;
		12'b011111010001: colour_data = 24'b000000000000000000000000;
		12'b011111010010: colour_data = 24'b000000000000000000000000;
		12'b011111010011: colour_data = 24'b111111110000000010010110;
		12'b011111010100: colour_data = 24'b111111110000000010010110;
		12'b011111010101: colour_data = 24'b111111110000000010010110;
		12'b011111010110: colour_data = 24'b111111110000000010010110;
		12'b011111010111: colour_data = 24'b010001000100010011101110;
		12'b011111011000: colour_data = 24'b010001000100010011101110;
		12'b011111011001: colour_data = 24'b011001100110011011101110;
		12'b011111011010: colour_data = 24'b111111110000000010010110;
		12'b011111011011: colour_data = 24'b111111001111110011111100;
		12'b011111011100: colour_data = 24'b111111110000000010010110;
		12'b011111011101: colour_data = 24'b111111110000000010010110;
		12'b011111011110: colour_data = 24'b111111001111110011111100;
		12'b011111011111: colour_data = 24'b111111000000000000000000;
		12'b011111100000: colour_data = 24'b111111000000000000000000;
		12'b011111100001: colour_data = 24'b111111000000000000000000;
		12'b011111100010: colour_data = 24'b111111000000000000000000;
		12'b011111100011: colour_data = 24'b000000000000000000000000;
		12'b011111100100: colour_data = 24'b111111110000000010010110;

		12'b100000000000: colour_data = 24'b111111110000000010010110;
		12'b100000000001: colour_data = 24'b111111110000000010010110;
		12'b100000000010: colour_data = 24'b111111110000000010010110;
		12'b100000000011: colour_data = 24'b111111110000000010010110;
		12'b100000000100: colour_data = 24'b111111110000000010010110;
		12'b100000000101: colour_data = 24'b111111110000000010010110;
		12'b100000000110: colour_data = 24'b111111110000000010010110;
		12'b100000000111: colour_data = 24'b000000000000000000000000;
		12'b100000001000: colour_data = 24'b100100000000000000000000;
		12'b100000001001: colour_data = 24'b100100000000000000000000;
		12'b100000001010: colour_data = 24'b000000000000000000000000;
		12'b100000001011: colour_data = 24'b100100000000000000000000;
		12'b100000001100: colour_data = 24'b100100000000000000000000;
		12'b100000001101: colour_data = 24'b000000000000000000000000;
		12'b100000001110: colour_data = 24'b101101001011010010110100;
		12'b100000001111: colour_data = 24'b001000100010001011001100;
		12'b100000010000: colour_data = 24'b001000100010001011001100;
		12'b100000010001: colour_data = 24'b000000000000000000000000;
		12'b100000010010: colour_data = 24'b111111110000000010010110;
		12'b100000010011: colour_data = 24'b111111110000000010010110;
		12'b100000010100: colour_data = 24'b111111110000000010010110;
		12'b100000010101: colour_data = 24'b111111110000000010010110;
		12'b100000010110: colour_data = 24'b111111110000000010010110;
		12'b100000010111: colour_data = 24'b111111110000000010010110;
		12'b100000011000: colour_data = 24'b111111110000000010010110;
		12'b100000011001: colour_data = 24'b010001000100010011101110;
		12'b100000011010: colour_data = 24'b010001000100010011101110;
		12'b100000011011: colour_data = 24'b111111001111110011111100;
		12'b100000011100: colour_data = 24'b111111001111110011111100;
		12'b100000011101: colour_data = 24'b101101001011010010110100;
		12'b100000011110: colour_data = 24'b111111001111110011111100;
		12'b100000011111: colour_data = 24'b111111001111110011111100;
		12'b100000100000: colour_data = 24'b111111001111110011111100;
		12'b100000100001: colour_data = 24'b111111000000000000000000;
		12'b100000100010: colour_data = 24'b000000000000000000000000;
		12'b100000100011: colour_data = 24'b111111110000000010010110;
		12'b100000100100: colour_data = 24'b111111110000000010010110;

		12'b100001000000: colour_data = 24'b111111110000000010010110;
		12'b100001000001: colour_data = 24'b111111110000000010010110;
		12'b100001000010: colour_data = 24'b111111110000000010010110;
		12'b100001000011: colour_data = 24'b111111110000000010010110;
		12'b100001000100: colour_data = 24'b111111110000000010010110;
		12'b100001000101: colour_data = 24'b111111110000000010010110;
		12'b100001000110: colour_data = 24'b111111110000000010010110;
		12'b100001000111: colour_data = 24'b000000000000000000000000;
		12'b100001001000: colour_data = 24'b100100000000000000000000;
		12'b100001001001: colour_data = 24'b000000000000000000000000;
		12'b100001001010: colour_data = 24'b100100000000000000000000;
		12'b100001001011: colour_data = 24'b100100000000000000000000;
		12'b100001001100: colour_data = 24'b100100000000000000000000;
		12'b100001001101: colour_data = 24'b100100001001000010010000;
		12'b100001001110: colour_data = 24'b100100001001000010010000;
		12'b100001001111: colour_data = 24'b001000100010001011001100;
		12'b100001010000: colour_data = 24'b000000000000000000000000;
		12'b100001010001: colour_data = 24'b111111110000000010010110;
		12'b100001010010: colour_data = 24'b111111110000000010010110;
		12'b100001010011: colour_data = 24'b111111110000000010010110;
		12'b100001010100: colour_data = 24'b111111110000000010010110;
		12'b100001010101: colour_data = 24'b111111110000000010010110;
		12'b100001010110: colour_data = 24'b111111110000000010010110;
		12'b100001010111: colour_data = 24'b111111110000000010010110;
		12'b100001011000: colour_data = 24'b111111110000000010010110;
		12'b100001011001: colour_data = 24'b111111110000000010010110;
		12'b100001011010: colour_data = 24'b111111001111110011111100;
		12'b100001011011: colour_data = 24'b111111001111110011111100;
		12'b100001011100: colour_data = 24'b111111001111110011111100;
		12'b100001011101: colour_data = 24'b111111000000000000000000;
		12'b100001011110: colour_data = 24'b111111000000000000000000;
		12'b100001011111: colour_data = 24'b111111000000000000000000;
		12'b100001100000: colour_data = 24'b111111001111110011111100;
		12'b100001100001: colour_data = 24'b111111001111110011111100;
		12'b100001100010: colour_data = 24'b000000000000000000000000;
		12'b100001100011: colour_data = 24'b111111110000000010010110;
		12'b100001100100: colour_data = 24'b111111110000000010010110;

		12'b100010000000: colour_data = 24'b111111110000000010010110;
		12'b100010000001: colour_data = 24'b111111110000000010010110;
		12'b100010000010: colour_data = 24'b111111110000000010010110;
		12'b100010000011: colour_data = 24'b111111110000000010010110;
		12'b100010000100: colour_data = 24'b111111110000000010010110;
		12'b100010000101: colour_data = 24'b111111110000000010010110;
		12'b100010000110: colour_data = 24'b111111110000000010010110;
		12'b100010000111: colour_data = 24'b000000000000000000000000;
		12'b100010001000: colour_data = 24'b100100000000000000000000;
		12'b100010001001: colour_data = 24'b000000000000000000000000;
		12'b100010001010: colour_data = 24'b100100000000000000000000;
		12'b100010001011: colour_data = 24'b100100000000000000000000;
		12'b100010001100: colour_data = 24'b000000000000000000000000;
		12'b100010001101: colour_data = 24'b100100001001000010010000;
		12'b100010001110: colour_data = 24'b000000000000000000000000;
		12'b100010001111: colour_data = 24'b000000000000000000000000;
		12'b100010010000: colour_data = 24'b111111110000000010010110;
		12'b100010010001: colour_data = 24'b111111110000000010010110;
		12'b100010010010: colour_data = 24'b111111110000000010010110;
		12'b100010010011: colour_data = 24'b111111110000000010010110;
		12'b100010010100: colour_data = 24'b111111110000000010010110;
		12'b100010010101: colour_data = 24'b111111110000000010010110;
		12'b100010010110: colour_data = 24'b111111110000000010010110;
		12'b100010010111: colour_data = 24'b111111110000000010010110;
		12'b100010011000: colour_data = 24'b111111110000000010010110;
		12'b100010011001: colour_data = 24'b101101001011010010110100;
		12'b100010011010: colour_data = 24'b111111001111110011111100;
		12'b100010011011: colour_data = 24'b111111001111110011111100;
		12'b100010011100: colour_data = 24'b111111001111110011111100;
		12'b100010011101: colour_data = 24'b111111000000000000000000;
		12'b100010011110: colour_data = 24'b111111000000000000000000;
		12'b100010011111: colour_data = 24'b111111000000000000000000;
		12'b100010100000: colour_data = 24'b101101001011010010110100;
		12'b100010100001: colour_data = 24'b000000000000000000000000;
		12'b100010100010: colour_data = 24'b111111110000000010010110;
		12'b100010100011: colour_data = 24'b111111110000000010010110;
		12'b100010100100: colour_data = 24'b111111110000000010010110;

		12'b100011000000: colour_data = 24'b111111110000000010010110;
		12'b100011000001: colour_data = 24'b111111110000000010010110;
		12'b100011000010: colour_data = 24'b111111110000000010010110;
		12'b100011000011: colour_data = 24'b111111110000000010010110;
		12'b100011000100: colour_data = 24'b111111110000000010010110;
		12'b100011000101: colour_data = 24'b111111110000000010010110;
		12'b100011000110: colour_data = 24'b000000000000000000000000;
		12'b100011000111: colour_data = 24'b100100000000000000000000;
		12'b100011001000: colour_data = 24'b100100000000000000000000;
		12'b100011001001: colour_data = 24'b000000000000000000000000;
		12'b100011001010: colour_data = 24'b100100000000000000000000;
		12'b100011001011: colour_data = 24'b100100000000000000000000;
		12'b100011001100: colour_data = 24'b000000000000000000000000;
		12'b100011001101: colour_data = 24'b000000000000000000000000;
		12'b100011001110: colour_data = 24'b111111110000000010010110;
		12'b100011001111: colour_data = 24'b111111110000000010010110;
		12'b100011010000: colour_data = 24'b111111110000000010010110;
		12'b100011010001: colour_data = 24'b111111110000000010010110;
		12'b100011010010: colour_data = 24'b111111110000000010010110;
		12'b100011010011: colour_data = 24'b111111110000000010010110;
		12'b100011010100: colour_data = 24'b111111110000000010010110;
		12'b100011010101: colour_data = 24'b111111110000000010010110;
		12'b100011010110: colour_data = 24'b111111110000000010010110;
		12'b100011010111: colour_data = 24'b111111110000000010010110;
		12'b100011011000: colour_data = 24'b111111110000000010010110;
		12'b100011011001: colour_data = 24'b111111110000000010010110;
		12'b100011011010: colour_data = 24'b101101001011010010110100;
		12'b100011011011: colour_data = 24'b111111001111110011111100;
		12'b100011011100: colour_data = 24'b111111000000000000000000;
		12'b100011011101: colour_data = 24'b111111000000000000000000;
		12'b100011011110: colour_data = 24'b111111000000000000000000;
		12'b100011011111: colour_data = 24'b111111000000000000000000;
		12'b100011100000: colour_data = 24'b000000000000000000000000;
		12'b100011100001: colour_data = 24'b111111110000000010010110;
		12'b100011100010: colour_data = 24'b111111110000000010010110;
		12'b100011100011: colour_data = 24'b111111110000000010010110;
		12'b100011100100: colour_data = 24'b111111110000000010010110;

		12'b100100000000: colour_data = 24'b111111110000000010010110;
		12'b100100000001: colour_data = 24'b111111110000000010010110;
		12'b100100000010: colour_data = 24'b111111110000000010010110;
		12'b100100000011: colour_data = 24'b111111110000000010010110;
		12'b100100000100: colour_data = 24'b111111110000000010010110;
		12'b100100000101: colour_data = 24'b111111110000000010010110;
		12'b100100000110: colour_data = 24'b000000000000000000000000;
		12'b100100000111: colour_data = 24'b100100000000000000000000;
		12'b100100001000: colour_data = 24'b000000000000000000000000;
		12'b100100001001: colour_data = 24'b111111001111110011111100;
		12'b100100001010: colour_data = 24'b111111001111110011111100;
		12'b100100001011: colour_data = 24'b000000000000000000000000;
		12'b100100001100: colour_data = 24'b111111110000000010010110;
		12'b100100001101: colour_data = 24'b111111110000000010010110;
		12'b100100001110: colour_data = 24'b111111110000000010010110;
		12'b100100001111: colour_data = 24'b111111110000000010010110;
		12'b100100010000: colour_data = 24'b111111110000000010010110;
		12'b100100010001: colour_data = 24'b111111110000000010010110;
		12'b100100010010: colour_data = 24'b111111110000000010010110;
		12'b100100010011: colour_data = 24'b111111110000000010010110;
		12'b100100010100: colour_data = 24'b111111110000000010010110;
		12'b100100010101: colour_data = 24'b111111110000000010010110;
		12'b100100010110: colour_data = 24'b111111110000000010010110;
		12'b100100010111: colour_data = 24'b111111110000000010010110;
		12'b100100011000: colour_data = 24'b111111110000000010010110;
		12'b100100011001: colour_data = 24'b111111110000000010010110;
		12'b100100011010: colour_data = 24'b000000000000000000000000;
		12'b100100011011: colour_data = 24'b111111000000000000000000;
		12'b100100011100: colour_data = 24'b111111000000000000000000;
		12'b100100011101: colour_data = 24'b111111000000000000000000;
		12'b100100011110: colour_data = 24'b111111000000000000000000;
		12'b100100011111: colour_data = 24'b111111000000000000000000;
		12'b100100100000: colour_data = 24'b000000000000000000000000;
		12'b100100100001: colour_data = 24'b111111110000000010010110;
		12'b100100100010: colour_data = 24'b111111110000000010010110;
		12'b100100100011: colour_data = 24'b111111110000000010010110;
		12'b100100100100: colour_data = 24'b111111110000000010010110;

		12'b100101000000: colour_data = 24'b111111110000000010010110;
		12'b100101000001: colour_data = 24'b111111110000000010010110;
		12'b100101000010: colour_data = 24'b111111110000000010010110;
		12'b100101000011: colour_data = 24'b111111110000000010010110;
		12'b100101000100: colour_data = 24'b111111110000000010010110;
		12'b100101000101: colour_data = 24'b111111110000000010010110;
		12'b100101000110: colour_data = 24'b000000000000000000000000;
		12'b100101000111: colour_data = 24'b100100000000000000000000;
		12'b100101001000: colour_data = 24'b000000000000000000000000;
		12'b100101001001: colour_data = 24'b111111001111110011111100;
		12'b100101001010: colour_data = 24'b111111001111110011111100;
		12'b100101001011: colour_data = 24'b000000000000000000000000;
		12'b100101001100: colour_data = 24'b111111110000000010010110;
		12'b100101001101: colour_data = 24'b111111110000000010010110;
		12'b100101001110: colour_data = 24'b111111110000000010010110;
		12'b100101001111: colour_data = 24'b111111110000000010010110;
		12'b100101010000: colour_data = 24'b111111110000000010010110;
		12'b100101010001: colour_data = 24'b111111110000000010010110;
		12'b100101010010: colour_data = 24'b111111110000000010010110;
		12'b100101010011: colour_data = 24'b111111110000000010010110;
		12'b100101010100: colour_data = 24'b111111110000000010010110;
		12'b100101010101: colour_data = 24'b111111110000000010010110;
		12'b100101010110: colour_data = 24'b111111110000000010010110;
		12'b100101010111: colour_data = 24'b111111110000000010010110;
		12'b100101011000: colour_data = 24'b111111110000000010010110;
		12'b100101011001: colour_data = 24'b111111110000000010010110;
		12'b100101011010: colour_data = 24'b000000000000000000000000;
		12'b100101011011: colour_data = 24'b111111000000000000000000;
		12'b100101011100: colour_data = 24'b111111000000000000000000;
		12'b100101011101: colour_data = 24'b111111000000000000000000;
		12'b100101011110: colour_data = 24'b111111000000000000000000;
		12'b100101011111: colour_data = 24'b000000000000000000000000;
		12'b100101100000: colour_data = 24'b111111110000000010010110;
		12'b100101100001: colour_data = 24'b111111110000000010010110;
		12'b100101100010: colour_data = 24'b111111110000000010010110;
		12'b100101100011: colour_data = 24'b111111110000000010010110;
		12'b100101100100: colour_data = 24'b111111110000000010010110;

		12'b100110000000: colour_data = 24'b111111110000000010010110;
		12'b100110000001: colour_data = 24'b111111110000000010010110;
		12'b100110000010: colour_data = 24'b111111110000000010010110;
		12'b100110000011: colour_data = 24'b111111110000000010010110;
		12'b100110000100: colour_data = 24'b111111110000000010010110;
		12'b100110000101: colour_data = 24'b000000000000000000000000;
		12'b100110000110: colour_data = 24'b100100000000000000000000;
		12'b100110000111: colour_data = 24'b000000000000000000000000;
		12'b100110001000: colour_data = 24'b100100000000000000000000;
		12'b100110001001: colour_data = 24'b100100000000000000000000;
		12'b100110001010: colour_data = 24'b000000000000000000000000;
		12'b100110001011: colour_data = 24'b111111110000000010010110;
		12'b100110001100: colour_data = 24'b111111110000000010010110;
		12'b100110001101: colour_data = 24'b111111110000000010010110;
		12'b100110001110: colour_data = 24'b111111110000000010010110;
		12'b100110001111: colour_data = 24'b111111110000000010010110;
		12'b100110010000: colour_data = 24'b111111110000000010010110;
		12'b100110010001: colour_data = 24'b111111110000000010010110;
		12'b100110010010: colour_data = 24'b111111110000000010010110;
		12'b100110010011: colour_data = 24'b111111110000000010010110;
		12'b100110010100: colour_data = 24'b111111110000000010010110;
		12'b100110010101: colour_data = 24'b111111110000000010010110;
		12'b100110010110: colour_data = 24'b111111110000000010010110;
		12'b100110010111: colour_data = 24'b111111110000000010010110;
		12'b100110011000: colour_data = 24'b111111110000000010010110;
		12'b100110011001: colour_data = 24'b111111110000000010010110;
		12'b100110011010: colour_data = 24'b111111110000000010010110;
		12'b100110011011: colour_data = 24'b000000000000000000000000;
		12'b100110011100: colour_data = 24'b111111000000000000000000;
		12'b100110011101: colour_data = 24'b111111000000000000000000;
		12'b100110011110: colour_data = 24'b000000000000000000000000;
		12'b100110011111: colour_data = 24'b111111110000000010010110;
		12'b100110100000: colour_data = 24'b111111110000000010010110;
		12'b100110100001: colour_data = 24'b111111110000000010010110;
		12'b100110100010: colour_data = 24'b111111110000000010010110;
		12'b100110100011: colour_data = 24'b111111110000000010010110;
		12'b100110100100: colour_data = 24'b111111110000000010010110;

		12'b100111000000: colour_data = 24'b111111110000000010010110;
		12'b100111000001: colour_data = 24'b111111110000000010010110;
		12'b100111000010: colour_data = 24'b111111110000000010010110;
		12'b100111000011: colour_data = 24'b111111110000000010010110;
		12'b100111000100: colour_data = 24'b111111110000000010010110;
		12'b100111000101: colour_data = 24'b000000000000000000000000;
		12'b100111000110: colour_data = 24'b100100000000000000000000;
		12'b100111000111: colour_data = 24'b000000000000000000000000;
		12'b100111001000: colour_data = 24'b100100000000000000000000;
		12'b100111001001: colour_data = 24'b000000000000000000000000;
		12'b100111001010: colour_data = 24'b111111110000000010010110;
		12'b100111001011: colour_data = 24'b111111110000000010010110;
		12'b100111001100: colour_data = 24'b111111110000000010010110;
		12'b100111001101: colour_data = 24'b111111110000000010010110;
		12'b100111001110: colour_data = 24'b111111110000000010010110;
		12'b100111001111: colour_data = 24'b111111110000000010010110;
		12'b100111010000: colour_data = 24'b111111110000000010010110;
		12'b100111010001: colour_data = 24'b111111110000000010010110;
		12'b100111010010: colour_data = 24'b111111110000000010010110;
		12'b100111010011: colour_data = 24'b111111110000000010010110;
		12'b100111010100: colour_data = 24'b111111110000000010010110;
		12'b100111010101: colour_data = 24'b111111110000000010010110;
		12'b100111010110: colour_data = 24'b111111110000000010010110;
		12'b100111010111: colour_data = 24'b111111110000000010010110;
		12'b100111011000: colour_data = 24'b111111110000000010010110;
		12'b100111011001: colour_data = 24'b111111110000000010010110;
		12'b100111011010: colour_data = 24'b111111110000000010010110;
		12'b100111011011: colour_data = 24'b111111110000000010010110;
		12'b100111011100: colour_data = 24'b000000000000000000000000;
		12'b100111011101: colour_data = 24'b000000000000000000000000;
		12'b100111011110: colour_data = 24'b111111110000000010010110;
		12'b100111011111: colour_data = 24'b111111110000000010010110;
		12'b100111100000: colour_data = 24'b111111110000000010010110;
		12'b100111100001: colour_data = 24'b111111110000000010010110;
		12'b100111100010: colour_data = 24'b111111110000000010010110;
		12'b100111100011: colour_data = 24'b111111110000000010010110;
		12'b100111100100: colour_data = 24'b111111110000000010010110;

		12'b101000000000: colour_data = 24'b111111110000000010010110;
		12'b101000000001: colour_data = 24'b111111110000000010010110;
		12'b101000000010: colour_data = 24'b111111110000000010010110;
		12'b101000000011: colour_data = 24'b111111110000000010010110;
		12'b101000000100: colour_data = 24'b111111110000000010010110;
		12'b101000000101: colour_data = 24'b000000000000000000000000;
		12'b101000000110: colour_data = 24'b000000000000000000000000;
		12'b101000000111: colour_data = 24'b100100000000000000000000;
		12'b101000001000: colour_data = 24'b000000000000000000000000;
		12'b101000001001: colour_data = 24'b111111110000000010010110;
		12'b101000001010: colour_data = 24'b111111110000000010010110;
		12'b101000001011: colour_data = 24'b111111110000000010010110;
		12'b101000001100: colour_data = 24'b111111110000000010010110;
		12'b101000001101: colour_data = 24'b111111110000000010010110;
		12'b101000001110: colour_data = 24'b111111110000000010010110;
		12'b101000001111: colour_data = 24'b111111110000000010010110;
		12'b101000010000: colour_data = 24'b111111110000000010010110;
		12'b101000010001: colour_data = 24'b111111110000000010010110;
		12'b101000010010: colour_data = 24'b111111110000000010010110;
		12'b101000010011: colour_data = 24'b111111110000000010010110;
		12'b101000010100: colour_data = 24'b111111110000000010010110;
		12'b101000010101: colour_data = 24'b111111110000000010010110;
		12'b101000010110: colour_data = 24'b111111110000000010010110;
		12'b101000010111: colour_data = 24'b111111110000000010010110;
		12'b101000011000: colour_data = 24'b111111110000000010010110;
		12'b101000011001: colour_data = 24'b111111110000000010010110;
		12'b101000011010: colour_data = 24'b111111110000000010010110;
		12'b101000011011: colour_data = 24'b111111110000000010010110;
		12'b101000011100: colour_data = 24'b111111110000000010010110;
		12'b101000011101: colour_data = 24'b111111110000000010010110;
		12'b101000011110: colour_data = 24'b111111110000000010010110;
		12'b101000011111: colour_data = 24'b111111110000000010010110;
		12'b101000100000: colour_data = 24'b111111110000000010010110;
		12'b101000100001: colour_data = 24'b111111110000000010010110;
		12'b101000100010: colour_data = 24'b111111110000000010010110;
		12'b101000100011: colour_data = 24'b111111110000000010010110;
		12'b101000100100: colour_data = 24'b111111110000000010010110;

		12'b101001000000: colour_data = 24'b111111110000000010010110;
		12'b101001000001: colour_data = 24'b111111110000000010010110;
		12'b101001000010: colour_data = 24'b111111110000000010010110;
		12'b101001000011: colour_data = 24'b111111110000000010010110;
		12'b101001000100: colour_data = 24'b111111110000000010010110;
		12'b101001000101: colour_data = 24'b000000000000000000000000;
		12'b101001000110: colour_data = 24'b000000000000000000000000;
		12'b101001000111: colour_data = 24'b000000000000000000000000;
		12'b101001001000: colour_data = 24'b111111110000000010010110;
		12'b101001001001: colour_data = 24'b111111110000000010010110;
		12'b101001001010: colour_data = 24'b111111110000000010010110;
		12'b101001001011: colour_data = 24'b111111110000000010010110;
		12'b101001001100: colour_data = 24'b111111110000000010010110;
		12'b101001001101: colour_data = 24'b111111110000000010010110;
		12'b101001001110: colour_data = 24'b111111110000000010010110;
		12'b101001001111: colour_data = 24'b111111110000000010010110;
		12'b101001010000: colour_data = 24'b111111110000000010010110;
		12'b101001010001: colour_data = 24'b111111110000000010010110;
		12'b101001010010: colour_data = 24'b111111110000000010010110;
		12'b101001010011: colour_data = 24'b111111110000000010010110;
		12'b101001010100: colour_data = 24'b111111110000000010010110;
		12'b101001010101: colour_data = 24'b111111110000000010010110;
		12'b101001010110: colour_data = 24'b111111110000000010010110;
		12'b101001010111: colour_data = 24'b111111110000000010010110;
		12'b101001011000: colour_data = 24'b111111110000000010010110;
		12'b101001011001: colour_data = 24'b111111110000000010010110;
		12'b101001011010: colour_data = 24'b111111110000000010010110;
		12'b101001011011: colour_data = 24'b111111110000000010010110;
		12'b101001011100: colour_data = 24'b111111110000000010010110;
		12'b101001011101: colour_data = 24'b111111110000000010010110;
		12'b101001011110: colour_data = 24'b111111110000000010010110;
		12'b101001011111: colour_data = 24'b111111110000000010010110;
		12'b101001100000: colour_data = 24'b111111110000000010010110;
		12'b101001100001: colour_data = 24'b111111110000000010010110;
		12'b101001100010: colour_data = 24'b111111110000000010010110;
		12'b101001100011: colour_data = 24'b111111110000000010010110;
		12'b101001100100: colour_data = 24'b111111110000000010010110;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule