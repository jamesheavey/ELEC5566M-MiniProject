module pause_rom
	(
		input wire clk,
		input wire [3:0] row,
		input wire [3:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [3:0] row_reg;
	reg [3:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		8'b00000000: colour_data = 24'b010101010011000000000000;
		8'b00000001: colour_data = 24'b010101010011000000000000;
		8'b00000010: colour_data = 24'b010101010011000000000000;
		8'b00000011: colour_data = 24'b010101010011000000000000;
		8'b00000100: colour_data = 24'b010101010011000000000000;
		8'b00000101: colour_data = 24'b010101010011000000000000;
		8'b00000110: colour_data = 24'b010101010011000000000000;
		8'b00000111: colour_data = 24'b010101010011000000000000;
		8'b00001000: colour_data = 24'b010101010011000000000000;
		8'b00001001: colour_data = 24'b010101010011000000000000;
		8'b00001010: colour_data = 24'b010101010011000000000000;
		8'b00001011: colour_data = 24'b010101010011000000000000;
		8'b00001100: colour_data = 24'b010101010011000000000000;

		8'b00010000: colour_data = 24'b010101010011000000000000;
		8'b00010001: colour_data = 24'b111111011111111011111101;
		8'b00010010: colour_data = 24'b111111011111111011111101;
		8'b00010011: colour_data = 24'b111111011111111011111101;
		8'b00010100: colour_data = 24'b111111011111111011111101;
		8'b00010101: colour_data = 24'b111111011111111011111101;
		8'b00010110: colour_data = 24'b111111011111111011111101;
		8'b00010111: colour_data = 24'b111111011111111011111101;
		8'b00011000: colour_data = 24'b111111011111111011111101;
		8'b00011001: colour_data = 24'b111111011111111011111101;
		8'b00011010: colour_data = 24'b111111011111111011111101;
		8'b00011011: colour_data = 24'b111111011111111011111101;
		8'b00011100: colour_data = 24'b010101010011000000000000;

		8'b00100000: colour_data = 24'b010101010011000000000000;
		8'b00100001: colour_data = 24'b111111011111111011111101;
		8'b00100010: colour_data = 24'b111010000110000100000000;
		8'b00100011: colour_data = 24'b111010000110000100000000;
		8'b00100100: colour_data = 24'b111010000110000100000000;
		8'b00100101: colour_data = 24'b111010000110000100000000;
		8'b00100110: colour_data = 24'b111010000110000100000000;
		8'b00100111: colour_data = 24'b111010000110000100000000;
		8'b00101000: colour_data = 24'b111010000110000100000000;
		8'b00101001: colour_data = 24'b111010000110000100000000;
		8'b00101010: colour_data = 24'b111010000110000100000000;
		8'b00101011: colour_data = 24'b111111011111111011111101;
		8'b00101100: colour_data = 24'b010101010011000000000000;

		8'b00110000: colour_data = 24'b010101010011000000000000;
		8'b00110001: colour_data = 24'b111111011111111011111101;
		8'b00110010: colour_data = 24'b111010000110000100000000;
		8'b00110011: colour_data = 24'b111010000110000100000000;
		8'b00110100: colour_data = 24'b111010000110000100000000;
		8'b00110101: colour_data = 24'b111010000110000100000000;
		8'b00110110: colour_data = 24'b111010000110000100000000;
		8'b00110111: colour_data = 24'b111010000110000100000000;
		8'b00111000: colour_data = 24'b111010000110000100000000;
		8'b00111001: colour_data = 24'b111010000110000100000000;
		8'b00111010: colour_data = 24'b111010000110000100000000;
		8'b00111011: colour_data = 24'b111111011111111011111101;
		8'b00111100: colour_data = 24'b010101010011000000000000;

		8'b01000000: colour_data = 24'b010101010011000000000000;
		8'b01000001: colour_data = 24'b111111011111111011111101;
		8'b01000010: colour_data = 24'b111010000110000100000000;
		8'b01000011: colour_data = 24'b111010000110000100000000;
		8'b01000100: colour_data = 24'b111111011111111011111101;
		8'b01000101: colour_data = 24'b111111011111111011111101;
		8'b01000110: colour_data = 24'b111010000110000100000000;
		8'b01000111: colour_data = 24'b111111011111111011111101;
		8'b01001000: colour_data = 24'b111111011111111011111101;
		8'b01001001: colour_data = 24'b111010000110000100000000;
		8'b01001010: colour_data = 24'b111010000110000100000000;
		8'b01001011: colour_data = 24'b111111011111111011111101;
		8'b01001100: colour_data = 24'b010101010011000000000000;

		8'b01010000: colour_data = 24'b010101010011000000000000;
		8'b01010001: colour_data = 24'b111111011111111011111101;
		8'b01010010: colour_data = 24'b111010000110000100000000;
		8'b01010011: colour_data = 24'b111010000110000100000000;
		8'b01010100: colour_data = 24'b111111011111111011111101;
		8'b01010101: colour_data = 24'b111111011111111011111101;
		8'b01010110: colour_data = 24'b111010000110000100000000;
		8'b01010111: colour_data = 24'b111111011111111011111101;
		8'b01011000: colour_data = 24'b111111011111111011111101;
		8'b01011001: colour_data = 24'b111010000110000100000000;
		8'b01011010: colour_data = 24'b111010000110000100000000;
		8'b01011011: colour_data = 24'b111111011111111011111101;
		8'b01011100: colour_data = 24'b010101010011000000000000;

		8'b01100000: colour_data = 24'b010101010011000000000000;
		8'b01100001: colour_data = 24'b111111011111111011111101;
		8'b01100010: colour_data = 24'b111010000110000100000000;
		8'b01100011: colour_data = 24'b111010000110000100000000;
		8'b01100100: colour_data = 24'b111111011111111011111101;
		8'b01100101: colour_data = 24'b111111011111111011111101;
		8'b01100110: colour_data = 24'b111010000110000100000000;
		8'b01100111: colour_data = 24'b111111011111111011111101;
		8'b01101000: colour_data = 24'b111111011111111011111101;
		8'b01101001: colour_data = 24'b111010000110000100000000;
		8'b01101010: colour_data = 24'b111010000110000100000000;
		8'b01101011: colour_data = 24'b111111011111111011111101;
		8'b01101100: colour_data = 24'b010101010011000000000000;

		8'b01110000: colour_data = 24'b010101010011000000000000;
		8'b01110001: colour_data = 24'b111111011111111011111101;
		8'b01110010: colour_data = 24'b111010000110000100000000;
		8'b01110011: colour_data = 24'b111010000110000100000000;
		8'b01110100: colour_data = 24'b111111011111111011111101;
		8'b01110101: colour_data = 24'b111111011111111011111101;
		8'b01110110: colour_data = 24'b111010000110000100000000;
		8'b01110111: colour_data = 24'b111111011111111011111101;
		8'b01111000: colour_data = 24'b111111011111111011111101;
		8'b01111001: colour_data = 24'b111010000110000100000000;
		8'b01111010: colour_data = 24'b111010000110000100000000;
		8'b01111011: colour_data = 24'b111111011111111011111101;
		8'b01111100: colour_data = 24'b010101010011000000000000;

		8'b10000000: colour_data = 24'b010101010011000000000000;
		8'b10000001: colour_data = 24'b111111011111111011111101;
		8'b10000010: colour_data = 24'b111010000110000100000000;
		8'b10000011: colour_data = 24'b111010000110000100000000;
		8'b10000100: colour_data = 24'b111111011111111011111101;
		8'b10000101: colour_data = 24'b111111011111111011111101;
		8'b10000110: colour_data = 24'b111010000110000100000000;
		8'b10000111: colour_data = 24'b111111011111111011111101;
		8'b10001000: colour_data = 24'b111111011111111011111101;
		8'b10001001: colour_data = 24'b111010000110000100000000;
		8'b10001010: colour_data = 24'b111010000110000100000000;
		8'b10001011: colour_data = 24'b111111011111111011111101;
		8'b10001100: colour_data = 24'b010101010011000000000000;

		8'b10010000: colour_data = 24'b010101010011000000000000;
		8'b10010001: colour_data = 24'b111111011111111011111101;
		8'b10010010: colour_data = 24'b111010000110000100000000;
		8'b10010011: colour_data = 24'b111010000110000100000000;
		8'b10010100: colour_data = 24'b101111110100111000000001;
		8'b10010101: colour_data = 24'b101111110100111000000001;
		8'b10010110: colour_data = 24'b111010000110000100000000;
		8'b10010111: colour_data = 24'b101111110100111000000001;
		8'b10011000: colour_data = 24'b101111110100111000000001;
		8'b10011001: colour_data = 24'b111010000110000100000000;
		8'b10011010: colour_data = 24'b111010000110000100000000;
		8'b10011011: colour_data = 24'b111111011111111011111101;
		8'b10011100: colour_data = 24'b010101010011000000000000;

		8'b10100000: colour_data = 24'b010101010011000000000000;
		8'b10100001: colour_data = 24'b111111011111111011111101;
		8'b10100010: colour_data = 24'b111010000110000100000000;
		8'b10100011: colour_data = 24'b111010000110000100000000;
		8'b10100100: colour_data = 24'b111010000110000100000000;
		8'b10100101: colour_data = 24'b111010000110000100000000;
		8'b10100110: colour_data = 24'b111010000110000100000000;
		8'b10100111: colour_data = 24'b111010000110000100000000;
		8'b10101000: colour_data = 24'b111010000110000100000000;
		8'b10101001: colour_data = 24'b111010000110000100000000;
		8'b10101010: colour_data = 24'b111010000110000100000000;
		8'b10101011: colour_data = 24'b111111011111111011111101;
		8'b10101100: colour_data = 24'b010101010011000000000000;

		8'b10110000: colour_data = 24'b010101010011000000000000;
		8'b10110001: colour_data = 24'b111111011111111011111101;
		8'b10110010: colour_data = 24'b111111011111111011111101;
		8'b10110011: colour_data = 24'b111111011111111011111101;
		8'b10110100: colour_data = 24'b111111011111111011111101;
		8'b10110101: colour_data = 24'b111111011111111011111101;
		8'b10110110: colour_data = 24'b111111011111111011111101;
		8'b10110111: colour_data = 24'b111111011111111011111101;
		8'b10111000: colour_data = 24'b111111011111111011111101;
		8'b10111001: colour_data = 24'b111111011111111011111101;
		8'b10111010: colour_data = 24'b111111011111111011111101;
		8'b10111011: colour_data = 24'b111111011111111011111101;
		8'b10111100: colour_data = 24'b010101010011000000000000;

		8'b11000000: colour_data = 24'b010101010011000000000000;
		8'b11000001: colour_data = 24'b010101010011000000000000;
		8'b11000010: colour_data = 24'b010101010011000000000000;
		8'b11000011: colour_data = 24'b010101010011000000000000;
		8'b11000100: colour_data = 24'b010101010011000000000000;
		8'b11000101: colour_data = 24'b010101010011000000000000;
		8'b11000110: colour_data = 24'b010101010011000000000000;
		8'b11000111: colour_data = 24'b010101010011000000000000;
		8'b11001000: colour_data = 24'b010101010011000000000000;
		8'b11001001: colour_data = 24'b010101010011000000000000;
		8'b11001010: colour_data = 24'b010101010011000000000000;
		8'b11001011: colour_data = 24'b010101010011000000000000;
		8'b11001100: colour_data = 24'b010101010011000000000000;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule