module bg_3_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [7:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		13'b0000000000000: colour_data = 24'b111111110000000010010110;
		13'b0000000000001: colour_data = 24'b011010101110001101011001;
		13'b0000000000010: colour_data = 24'b011010101110001101011001;
		13'b0000000000011: colour_data = 24'b001000011000111000100001;
		13'b0000000000100: colour_data = 24'b001000011000111000100001;
		13'b0000000000101: colour_data = 24'b011010101110001101011001;
		13'b0000000000110: colour_data = 24'b011010101110001101011001;
		13'b0000000000111: colour_data = 24'b001000011000111000100001;
		13'b0000000001000: colour_data = 24'b001000011000111000100001;
		13'b0000000001001: colour_data = 24'b001000011000111000100001;
		13'b0000000001010: colour_data = 24'b011010101110001101011001;
		13'b0000000001011: colour_data = 24'b011010101110001101011001;
		13'b0000000001100: colour_data = 24'b001000011000111000100001;
		13'b0000000001101: colour_data = 24'b001000011000111000100001;
		13'b0000000001110: colour_data = 24'b001000011000111000100001;
		13'b0000000001111: colour_data = 24'b011010101110001101011001;
		13'b0000000010000: colour_data = 24'b011010101110001101011001;
		13'b0000000010001: colour_data = 24'b001000011000111000100001;
		13'b0000000010010: colour_data = 24'b001000011000111000100001;
		13'b0000000010011: colour_data = 24'b011010101110001101011001;
		13'b0000000010100: colour_data = 24'b011010101110001101011001;
		13'b0000000010101: colour_data = 24'b011010101110001101011001;
		13'b0000000010110: colour_data = 24'b001000011000111000100001;
		13'b0000000010111: colour_data = 24'b001000011000111000100001;
		13'b0000000011000: colour_data = 24'b011010101110001101011001;
		13'b0000000011001: colour_data = 24'b011010101110001101011001;
		13'b0000000011010: colour_data = 24'b001000011000111000100001;
		13'b0000000011011: colour_data = 24'b001000011000111000100001;
		13'b0000000011100: colour_data = 24'b001000011000111000100001;
		13'b0000000011101: colour_data = 24'b011010101110001101011001;
		13'b0000000011110: colour_data = 24'b011010101110001101011001;
		13'b0000000011111: colour_data = 24'b001000011000111000100001;
		13'b0000000100000: colour_data = 24'b001000011000111000100001;
		13'b0000000100001: colour_data = 24'b011010101110001101011001;
		13'b0000000100010: colour_data = 24'b011010101110001101011001;
		13'b0000000100011: colour_data = 24'b011010101110001101011001;
		13'b0000000100100: colour_data = 24'b001000011000111000100001;
		13'b0000000100101: colour_data = 24'b001000011000111000100001;
		13'b0000000100110: colour_data = 24'b011010101110001101011001;
		13'b0000000100111: colour_data = 24'b011010101110001101011001;
		13'b0000000101000: colour_data = 24'b011010101110001101011001;
		13'b0000000101001: colour_data = 24'b001000011000111000100001;
		13'b0000000101010: colour_data = 24'b001000011000111000100001;
		13'b0000000101011: colour_data = 24'b011010101110001101011001;
		13'b0000000101100: colour_data = 24'b011010101110001101011001;
		13'b0000000101101: colour_data = 24'b001000011000111000100001;
		13'b0000000101110: colour_data = 24'b001000011000111000100001;
		13'b0000000101111: colour_data = 24'b001000011000111000100001;
		13'b0000000110000: colour_data = 24'b011010101110001101011001;
		13'b0000000110001: colour_data = 24'b011010101110001101011001;
		13'b0000000110010: colour_data = 24'b001000011000111000100001;
		13'b0000000110011: colour_data = 24'b001000011000111000100001;
		13'b0000000110100: colour_data = 24'b011010101110001101011001;
		13'b0000000110101: colour_data = 24'b011010101110001101011001;
		13'b0000000110110: colour_data = 24'b011010101110001101011001;
		13'b0000000110111: colour_data = 24'b001000011000111000100001;
		13'b0000000111000: colour_data = 24'b001000011000111000100001;
		13'b0000000111001: colour_data = 24'b011010101110001101011001;
		13'b0000000111010: colour_data = 24'b011010101110001101011001;
		13'b0000000111011: colour_data = 24'b011010101110001101011001;
		13'b0000000111100: colour_data = 24'b001000011000111000100001;
		13'b0000000111101: colour_data = 24'b001000011000111000100001;
		13'b0000000111110: colour_data = 24'b011010101110001101011001;
		13'b0000000111111: colour_data = 24'b011010101110001101011001;
		13'b0000001000000: colour_data = 24'b001000011000111000100001;
		13'b0000001000001: colour_data = 24'b001000011000111000100001;
		13'b0000001000010: colour_data = 24'b001000011000111000100001;
		13'b0000001000011: colour_data = 24'b011010101110001101011001;
		13'b0000001000100: colour_data = 24'b011010101110001101011001;
		13'b0000001000101: colour_data = 24'b001000011000111000100001;
		13'b0000001000110: colour_data = 24'b001000011000111000100001;
		13'b0000001000111: colour_data = 24'b011010101110001101011001;
		13'b0000001001000: colour_data = 24'b011010101110001101011001;
		13'b0000001001001: colour_data = 24'b011010101110001101011001;
		13'b0000001001010: colour_data = 24'b001000011000111000100001;
		13'b0000001001011: colour_data = 24'b001000011000111000100001;
		13'b0000001001100: colour_data = 24'b011010101110001101011001;
		13'b0000001001101: colour_data = 24'b011010101110001101011001;
		13'b0000001001110: colour_data = 24'b001000011000111000100001;
		13'b0000001001111: colour_data = 24'b001000011000111000100001;
		13'b0000001010000: colour_data = 24'b001000011000111000100001;
		13'b0000001010001: colour_data = 24'b011010101110001101011001;
		13'b0000001010010: colour_data = 24'b011010101110001101011001;
		13'b0000001010011: colour_data = 24'b001000011000111000100001;
		13'b0000001010100: colour_data = 24'b001000011000111000100001;
		13'b0000001010101: colour_data = 24'b001000011000111000100001;
		13'b0000001010110: colour_data = 24'b011010101110001101011001;
		13'b0000001010111: colour_data = 24'b011010101110001101011001;
		13'b0000001011000: colour_data = 24'b001000011000111000100001;
		13'b0000001011001: colour_data = 24'b001000011000111000100001;
		13'b0000001011010: colour_data = 24'b011010101110001101011001;
		13'b0000001011011: colour_data = 24'b011010101110001101011001;
		13'b0000001011100: colour_data = 24'b011010101110001101011001;
		13'b0000001011101: colour_data = 24'b001000011000111000100001;
		13'b0000001011110: colour_data = 24'b001000011000111000100001;
		13'b0000001011111: colour_data = 24'b011010101110001101011001;
		13'b0000001100000: colour_data = 24'b011010101110001101011001;
		13'b0000001100001: colour_data = 24'b001000011000111000100001;
		13'b0000001100010: colour_data = 24'b001000011000111000100001;
		13'b0000001100011: colour_data = 24'b001000011000111000100001;
		13'b0000001100100: colour_data = 24'b011010101110001101011001;
		13'b0000001100101: colour_data = 24'b011010101110001101011001;
		13'b0000001100110: colour_data = 24'b001000011000111000100001;
		13'b0000001100111: colour_data = 24'b001000011000111000100001;
		13'b0000001101000: colour_data = 24'b001000011000111000100001;
		13'b0000001101001: colour_data = 24'b011010101110001101011001;
		13'b0000001101010: colour_data = 24'b011010101110001101011001;
		13'b0000001101011: colour_data = 24'b001000011000111000100001;
		13'b0000001101100: colour_data = 24'b001000011000111000100001;
		13'b0000001101101: colour_data = 24'b011010101110001101011001;
		13'b0000001101110: colour_data = 24'b011010101110001101011001;
		13'b0000001101111: colour_data = 24'b011010101110001101011001;
		13'b0000001110000: colour_data = 24'b001000011000111000100001;
		13'b0000001110001: colour_data = 24'b001000011000111000100001;
		13'b0000001110010: colour_data = 24'b011010101110001101011001;
		13'b0000001110011: colour_data = 24'b011010101110001101011001;
		13'b0000001110100: colour_data = 24'b001000011000111000100001;
		13'b0000001110101: colour_data = 24'b001000011000111000100001;
		13'b0000001110110: colour_data = 24'b001000011000111000100001;
		13'b0000001110111: colour_data = 24'b011010101110001101011001;
		13'b0000001111000: colour_data = 24'b011010101110001101011001;
		13'b0000001111001: colour_data = 24'b001000011000111000100001;
		13'b0000001111010: colour_data = 24'b001000011000111000100001;
		13'b0000001111011: colour_data = 24'b011010101110001101011001;
		13'b0000001111100: colour_data = 24'b011010101110001101011001;
		13'b0000001111101: colour_data = 24'b011010101110001101011001;
		13'b0000001111110: colour_data = 24'b001000011000111000100001;
		13'b0000001111111: colour_data = 24'b001000011000111000100001;
		13'b0000010000000: colour_data = 24'b011010101110001101011001;
		13'b0000010000001: colour_data = 24'b011010101110001101011001;
		13'b0000010000010: colour_data = 24'b011010101110001101011001;
		13'b0000010000011: colour_data = 24'b001000011000111000100001;
		13'b0000010000100: colour_data = 24'b001000011000111000100001;
		13'b0000010000101: colour_data = 24'b011010101110001101011001;
		13'b0000010000110: colour_data = 24'b011010101110001101011001;
		13'b0000010000111: colour_data = 24'b001000011000111000100001;
		13'b0000010001000: colour_data = 24'b001000011000111000100001;
		13'b0000010001001: colour_data = 24'b000110000110110100011000;

		13'b0000100000000: colour_data = 24'b011010101110001101011001;
		13'b0000100000001: colour_data = 24'b101101011110111110110101;
		13'b0000100000010: colour_data = 24'b101101011110111110110101;
		13'b0000100000011: colour_data = 24'b011110001100011001101101;
		13'b0000100000100: colour_data = 24'b011110001100011001101101;
		13'b0000100000101: colour_data = 24'b101101011110111110110101;
		13'b0000100000110: colour_data = 24'b101101011110111110110101;
		13'b0000100000111: colour_data = 24'b011110001100011001101101;
		13'b0000100001000: colour_data = 24'b011110001100011001101101;
		13'b0000100001001: colour_data = 24'b011110001100011001101101;
		13'b0000100001010: colour_data = 24'b101101011110111110110101;
		13'b0000100001011: colour_data = 24'b101101011110111110110101;
		13'b0000100001100: colour_data = 24'b011110001100011001101101;
		13'b0000100001101: colour_data = 24'b011110001100011001101101;
		13'b0000100001110: colour_data = 24'b011110001100011001101101;
		13'b0000100001111: colour_data = 24'b101101011110111110110101;
		13'b0000100010000: colour_data = 24'b101101011110111110110101;
		13'b0000100010001: colour_data = 24'b011110001100011001101101;
		13'b0000100010010: colour_data = 24'b011110001100011001101101;
		13'b0000100010011: colour_data = 24'b101101011110111110110101;
		13'b0000100010100: colour_data = 24'b101101011110111110110101;
		13'b0000100010101: colour_data = 24'b101101011110111110110101;
		13'b0000100010110: colour_data = 24'b011110001100011001101101;
		13'b0000100010111: colour_data = 24'b011110001100011001101101;
		13'b0000100011000: colour_data = 24'b101101011110111110110101;
		13'b0000100011001: colour_data = 24'b101101011110111110110101;
		13'b0000100011010: colour_data = 24'b011110001100011001101101;
		13'b0000100011011: colour_data = 24'b011110001100011001101101;
		13'b0000100011100: colour_data = 24'b011110001100011001101101;
		13'b0000100011101: colour_data = 24'b101101011110111110110101;
		13'b0000100011110: colour_data = 24'b101101011110111110110101;
		13'b0000100011111: colour_data = 24'b011110001100011001101101;
		13'b0000100100000: colour_data = 24'b011110001100011001101101;
		13'b0000100100001: colour_data = 24'b101101011110111110110101;
		13'b0000100100010: colour_data = 24'b101101011110111110110101;
		13'b0000100100011: colour_data = 24'b101101011110111110110101;
		13'b0000100100100: colour_data = 24'b011110001100011001101101;
		13'b0000100100101: colour_data = 24'b011110001100011001101101;
		13'b0000100100110: colour_data = 24'b101101011110111110110101;
		13'b0000100100111: colour_data = 24'b101101011110111110110101;
		13'b0000100101000: colour_data = 24'b101101011110111110110101;
		13'b0000100101001: colour_data = 24'b011110001100011001101101;
		13'b0000100101010: colour_data = 24'b011110001100011001101101;
		13'b0000100101011: colour_data = 24'b101101011110111110110101;
		13'b0000100101100: colour_data = 24'b101101011110111110110101;
		13'b0000100101101: colour_data = 24'b011110001100011001101101;
		13'b0000100101110: colour_data = 24'b011110001100011001101101;
		13'b0000100101111: colour_data = 24'b011110001100011001101101;
		13'b0000100110000: colour_data = 24'b101101011110111110110101;
		13'b0000100110001: colour_data = 24'b101101011110111110110101;
		13'b0000100110010: colour_data = 24'b011110001100011001101101;
		13'b0000100110011: colour_data = 24'b011110001100011001101101;
		13'b0000100110100: colour_data = 24'b011010101110001101011001;
		13'b0000100110101: colour_data = 24'b101101011110111110110101;
		13'b0000100110110: colour_data = 24'b101101011110111110110101;
		13'b0000100110111: colour_data = 24'b011110001100011001101101;
		13'b0000100111000: colour_data = 24'b011110001100011001101101;
		13'b0000100111001: colour_data = 24'b101101011110111110110101;
		13'b0000100111010: colour_data = 24'b101101011110111110110101;
		13'b0000100111011: colour_data = 24'b101101011110111110110101;
		13'b0000100111100: colour_data = 24'b011110001100011001101101;
		13'b0000100111101: colour_data = 24'b011110001100011001101101;
		13'b0000100111110: colour_data = 24'b101101011110111110110101;
		13'b0000100111111: colour_data = 24'b101101011110111110110101;
		13'b0000101000000: colour_data = 24'b011110001100011001101101;
		13'b0000101000001: colour_data = 24'b011110001100011001101101;
		13'b0000101000010: colour_data = 24'b011110001100011001101101;
		13'b0000101000011: colour_data = 24'b101101011110111110110101;
		13'b0000101000100: colour_data = 24'b101101011110111110110101;
		13'b0000101000101: colour_data = 24'b011110001100011001101101;
		13'b0000101000110: colour_data = 24'b011110001100011001101101;
		13'b0000101000111: colour_data = 24'b101101011110111110110101;
		13'b0000101001000: colour_data = 24'b101101011110111110110101;
		13'b0000101001001: colour_data = 24'b101101011110111110110101;
		13'b0000101001010: colour_data = 24'b011110001100011001101101;
		13'b0000101001011: colour_data = 24'b011110001100011001101101;
		13'b0000101001100: colour_data = 24'b101101011110111110110101;
		13'b0000101001101: colour_data = 24'b101101011110111110110101;
		13'b0000101001110: colour_data = 24'b011110001100011001101101;
		13'b0000101001111: colour_data = 24'b011110001100011001101101;
		13'b0000101010000: colour_data = 24'b011110001100011001101101;
		13'b0000101010001: colour_data = 24'b101101011110111110110101;
		13'b0000101010010: colour_data = 24'b101101011110111110110101;
		13'b0000101010011: colour_data = 24'b011110001100011001101101;
		13'b0000101010100: colour_data = 24'b011110001100011001101101;
		13'b0000101010101: colour_data = 24'b011110001100011001101101;
		13'b0000101010110: colour_data = 24'b101101011110111110110101;
		13'b0000101010111: colour_data = 24'b101101011110111110110101;
		13'b0000101011000: colour_data = 24'b011110001100011001101101;
		13'b0000101011001: colour_data = 24'b011110001100011001101101;
		13'b0000101011010: colour_data = 24'b101101011110111110110101;
		13'b0000101011011: colour_data = 24'b101101011110111110110101;
		13'b0000101011100: colour_data = 24'b101101011110111110110101;
		13'b0000101011101: colour_data = 24'b011110001100011001101101;
		13'b0000101011110: colour_data = 24'b011110001100011001101101;
		13'b0000101011111: colour_data = 24'b101101011110111110110101;
		13'b0000101100000: colour_data = 24'b101101011110111110110101;
		13'b0000101100001: colour_data = 24'b011110001100011001101101;
		13'b0000101100010: colour_data = 24'b011110001100011001101101;
		13'b0000101100011: colour_data = 24'b011110001100011001101101;
		13'b0000101100100: colour_data = 24'b101101011110111110110101;
		13'b0000101100101: colour_data = 24'b101101011110111110110101;
		13'b0000101100110: colour_data = 24'b011110001100011001101101;
		13'b0000101100111: colour_data = 24'b011110001100011001101101;
		13'b0000101101000: colour_data = 24'b011110001100011001101101;
		13'b0000101101001: colour_data = 24'b101101011110111110110101;
		13'b0000101101010: colour_data = 24'b101101011110111110110101;
		13'b0000101101011: colour_data = 24'b011110001100011001101101;
		13'b0000101101100: colour_data = 24'b011110001100011001101101;
		13'b0000101101101: colour_data = 24'b101101011110111110110101;
		13'b0000101101110: colour_data = 24'b101101011110111110110101;
		13'b0000101101111: colour_data = 24'b101101011110111110110101;
		13'b0000101110000: colour_data = 24'b011110001100011001101101;
		13'b0000101110001: colour_data = 24'b011110001100011001101101;
		13'b0000101110010: colour_data = 24'b101101011110111110110101;
		13'b0000101110011: colour_data = 24'b101101011110111110110101;
		13'b0000101110100: colour_data = 24'b011110001100011001101101;
		13'b0000101110101: colour_data = 24'b011110001100011001101101;
		13'b0000101110110: colour_data = 24'b011110001100011001101101;
		13'b0000101110111: colour_data = 24'b101101011110111110110101;
		13'b0000101111000: colour_data = 24'b101101011110111110110101;
		13'b0000101111001: colour_data = 24'b011110001100011001101101;
		13'b0000101111010: colour_data = 24'b011110001100011001101101;
		13'b0000101111011: colour_data = 24'b101101011110111110110101;
		13'b0000101111100: colour_data = 24'b101101011110111110110101;
		13'b0000101111101: colour_data = 24'b101101011110111110110101;
		13'b0000101111110: colour_data = 24'b011110001100011001101101;
		13'b0000101111111: colour_data = 24'b011110001100011001101101;
		13'b0000110000000: colour_data = 24'b101101011110111110110101;
		13'b0000110000001: colour_data = 24'b101101011110111110110101;
		13'b0000110000010: colour_data = 24'b101101011110111110110101;
		13'b0000110000011: colour_data = 24'b011110001100011001101101;
		13'b0000110000100: colour_data = 24'b011110001100011001101101;
		13'b0000110000101: colour_data = 24'b101101011110111110110101;
		13'b0000110000110: colour_data = 24'b101101011110111110110101;
		13'b0000110000111: colour_data = 24'b011110001100011001101101;
		13'b0000110001000: colour_data = 24'b011110001100011001101101;
		13'b0000110001001: colour_data = 24'b001000011000111000100001;

		13'b0001000000000: colour_data = 24'b101101011110111110110101;
		13'b0001000000001: colour_data = 24'b111101111111111111101111;
		13'b0001000000010: colour_data = 24'b111101111111111111101111;
		13'b0001000000011: colour_data = 24'b101101011110111110110101;
		13'b0001000000100: colour_data = 24'b101101011110111110110101;
		13'b0001000000101: colour_data = 24'b111101111111111111101111;
		13'b0001000000110: colour_data = 24'b111101111111111111101111;
		13'b0001000000111: colour_data = 24'b101101011110111110110101;
		13'b0001000001000: colour_data = 24'b101101011110111110110101;
		13'b0001000001001: colour_data = 24'b101101011110111110110101;
		13'b0001000001010: colour_data = 24'b111101111111111111101111;
		13'b0001000001011: colour_data = 24'b111101111111111111101111;
		13'b0001000001100: colour_data = 24'b101101011110111110110101;
		13'b0001000001101: colour_data = 24'b101101011110111110110101;
		13'b0001000001110: colour_data = 24'b101101011110111110110101;
		13'b0001000001111: colour_data = 24'b111101111111111111101111;
		13'b0001000010000: colour_data = 24'b111101111111111111101111;
		13'b0001000010001: colour_data = 24'b101101011110111110110101;
		13'b0001000010010: colour_data = 24'b101101011110111110110101;
		13'b0001000010011: colour_data = 24'b111101111111111111101111;
		13'b0001000010100: colour_data = 24'b111101111111111111101111;
		13'b0001000010101: colour_data = 24'b111101111111111111101111;
		13'b0001000010110: colour_data = 24'b101101011110111110110101;
		13'b0001000010111: colour_data = 24'b101101011110111110110101;
		13'b0001000011000: colour_data = 24'b111101111111111111101111;
		13'b0001000011001: colour_data = 24'b111101111111111111101111;
		13'b0001000011010: colour_data = 24'b101101011110111110110101;
		13'b0001000011011: colour_data = 24'b101101011110111110110101;
		13'b0001000011100: colour_data = 24'b101101011110111110110101;
		13'b0001000011101: colour_data = 24'b111101111111111111101111;
		13'b0001000011110: colour_data = 24'b111101111111111111101111;
		13'b0001000011111: colour_data = 24'b101101011110111110110101;
		13'b0001000100000: colour_data = 24'b101101011110111110110101;
		13'b0001000100001: colour_data = 24'b111101111111111111101111;
		13'b0001000100010: colour_data = 24'b111101111111111111101111;
		13'b0001000100011: colour_data = 24'b111101111111111111101111;
		13'b0001000100100: colour_data = 24'b101101011110111110110101;
		13'b0001000100101: colour_data = 24'b101101011110111110110101;
		13'b0001000100110: colour_data = 24'b111101111111111111101111;
		13'b0001000100111: colour_data = 24'b111101111111111111101111;
		13'b0001000101000: colour_data = 24'b111101111111111111101111;
		13'b0001000101001: colour_data = 24'b101101011110111110110101;
		13'b0001000101010: colour_data = 24'b101101011110111110110101;
		13'b0001000101011: colour_data = 24'b111101111111111111101111;
		13'b0001000101100: colour_data = 24'b111101111111111111101111;
		13'b0001000101101: colour_data = 24'b101101011110111110110101;
		13'b0001000101110: colour_data = 24'b101101011110111110110101;
		13'b0001000101111: colour_data = 24'b101101011110111110110101;
		13'b0001000110000: colour_data = 24'b111101111111111111101111;
		13'b0001000110001: colour_data = 24'b111101111111111111101111;
		13'b0001000110010: colour_data = 24'b101101011110111110110101;
		13'b0001000110011: colour_data = 24'b101101011110111110110101;
		13'b0001000110100: colour_data = 24'b101101011110111110110101;
		13'b0001000110101: colour_data = 24'b111101111111111111101111;
		13'b0001000110110: colour_data = 24'b111101111111111111101111;
		13'b0001000110111: colour_data = 24'b101101011110111110110101;
		13'b0001000111000: colour_data = 24'b101101011110111110110101;
		13'b0001000111001: colour_data = 24'b111101111111111111101111;
		13'b0001000111010: colour_data = 24'b111101111111111111101111;
		13'b0001000111011: colour_data = 24'b111101111111111111101111;
		13'b0001000111100: colour_data = 24'b101101011110111110110101;
		13'b0001000111101: colour_data = 24'b101101011110111110110101;
		13'b0001000111110: colour_data = 24'b111101111111111111101111;
		13'b0001000111111: colour_data = 24'b111101111111111111101111;
		13'b0001001000000: colour_data = 24'b101101011110111110110101;
		13'b0001001000001: colour_data = 24'b101101011110111110110101;
		13'b0001001000010: colour_data = 24'b101101011110111110110101;
		13'b0001001000011: colour_data = 24'b111101111111111111101111;
		13'b0001001000100: colour_data = 24'b111101111111111111101111;
		13'b0001001000101: colour_data = 24'b101101011110111110110101;
		13'b0001001000110: colour_data = 24'b101101011110111110110101;
		13'b0001001000111: colour_data = 24'b111101111111111111101111;
		13'b0001001001000: colour_data = 24'b111101111111111111101111;
		13'b0001001001001: colour_data = 24'b111101111111111111101111;
		13'b0001001001010: colour_data = 24'b101101011110111110110101;
		13'b0001001001011: colour_data = 24'b101101011110111110110101;
		13'b0001001001100: colour_data = 24'b111101111111111111101111;
		13'b0001001001101: colour_data = 24'b111101111111111111101111;
		13'b0001001001110: colour_data = 24'b101101011110111110110101;
		13'b0001001001111: colour_data = 24'b101101011110111110110101;
		13'b0001001010000: colour_data = 24'b101101011110111110110101;
		13'b0001001010001: colour_data = 24'b111101111111111111101111;
		13'b0001001010010: colour_data = 24'b111101111111111111101111;
		13'b0001001010011: colour_data = 24'b101101011110111110110101;
		13'b0001001010100: colour_data = 24'b101101011110111110110101;
		13'b0001001010101: colour_data = 24'b101101011110111110110101;
		13'b0001001010110: colour_data = 24'b111101111111111111101111;
		13'b0001001010111: colour_data = 24'b111101111111111111101111;
		13'b0001001011000: colour_data = 24'b101101011110111110110101;
		13'b0001001011001: colour_data = 24'b101101011110111110110101;
		13'b0001001011010: colour_data = 24'b111101111111111111101111;
		13'b0001001011011: colour_data = 24'b111101111111111111101111;
		13'b0001001011100: colour_data = 24'b111101111111111111101111;
		13'b0001001011101: colour_data = 24'b101101011110111110110101;
		13'b0001001011110: colour_data = 24'b101101011110111110110101;
		13'b0001001011111: colour_data = 24'b111101111111111111101111;
		13'b0001001100000: colour_data = 24'b111101111111111111101111;
		13'b0001001100001: colour_data = 24'b101101011110111110110101;
		13'b0001001100010: colour_data = 24'b101101011110111110110101;
		13'b0001001100011: colour_data = 24'b101101011110111110110101;
		13'b0001001100100: colour_data = 24'b111101111111111111101111;
		13'b0001001100101: colour_data = 24'b111101111111111111101111;
		13'b0001001100110: colour_data = 24'b101101011110111110110101;
		13'b0001001100111: colour_data = 24'b101101011110111110110101;
		13'b0001001101000: colour_data = 24'b101101011110111110110101;
		13'b0001001101001: colour_data = 24'b111101111111111111101111;
		13'b0001001101010: colour_data = 24'b111101111111111111101111;
		13'b0001001101011: colour_data = 24'b101101011110111110110101;
		13'b0001001101100: colour_data = 24'b101101011110111110110101;
		13'b0001001101101: colour_data = 24'b111101111111111111101111;
		13'b0001001101110: colour_data = 24'b111101111111111111101111;
		13'b0001001101111: colour_data = 24'b111101111111111111101111;
		13'b0001001110000: colour_data = 24'b101101011110111110110101;
		13'b0001001110001: colour_data = 24'b101101011110111110110101;
		13'b0001001110010: colour_data = 24'b111101111111111111101111;
		13'b0001001110011: colour_data = 24'b111101111111111111101111;
		13'b0001001110100: colour_data = 24'b101101011110111110110101;
		13'b0001001110101: colour_data = 24'b101101011110111110110101;
		13'b0001001110110: colour_data = 24'b101101011110111110110101;
		13'b0001001110111: colour_data = 24'b111101111111111111101111;
		13'b0001001111000: colour_data = 24'b111101111111111111101111;
		13'b0001001111001: colour_data = 24'b101101011110111110110101;
		13'b0001001111010: colour_data = 24'b101101011110111110110101;
		13'b0001001111011: colour_data = 24'b111101111111111111101111;
		13'b0001001111100: colour_data = 24'b111101111111111111101111;
		13'b0001001111101: colour_data = 24'b111101111111111111101111;
		13'b0001001111110: colour_data = 24'b101101011110111110110101;
		13'b0001001111111: colour_data = 24'b101101011110111110110101;
		13'b0001010000000: colour_data = 24'b111101111111111111101111;
		13'b0001010000001: colour_data = 24'b111101111111111111101111;
		13'b0001010000010: colour_data = 24'b111101111111111111101111;
		13'b0001010000011: colour_data = 24'b101101011110111110110101;
		13'b0001010000100: colour_data = 24'b101101011110111110110101;
		13'b0001010000101: colour_data = 24'b111101111111111111101111;
		13'b0001010000110: colour_data = 24'b111101111111111111101111;
		13'b0001010000111: colour_data = 24'b101101011110111110110101;
		13'b0001010001000: colour_data = 24'b101101011110111110110101;
		13'b0001010001001: colour_data = 24'b011110001100011001101101;

		13'b0001100000000: colour_data = 24'b011010101110001101011001;
		13'b0001100000001: colour_data = 24'b101101011110111110110101;
		13'b0001100000010: colour_data = 24'b101101011110111110110101;
		13'b0001100000011: colour_data = 24'b011110001100011001101101;
		13'b0001100000100: colour_data = 24'b011110001100011001101101;
		13'b0001100000101: colour_data = 24'b101101011110111110110101;
		13'b0001100000110: colour_data = 24'b101101011110111110110101;
		13'b0001100000111: colour_data = 24'b011110001100011001101101;
		13'b0001100001000: colour_data = 24'b011110001100011001101101;
		13'b0001100001001: colour_data = 24'b011110001100011001101101;
		13'b0001100001010: colour_data = 24'b101101011110111110110101;
		13'b0001100001011: colour_data = 24'b101101011110111110110101;
		13'b0001100001100: colour_data = 24'b011110001100011001101101;
		13'b0001100001101: colour_data = 24'b011110001100011001101101;
		13'b0001100001110: colour_data = 24'b011110001100011001101101;
		13'b0001100001111: colour_data = 24'b101101011110111110110101;
		13'b0001100010000: colour_data = 24'b101101011110111110110101;
		13'b0001100010001: colour_data = 24'b011110001100011001101101;
		13'b0001100010010: colour_data = 24'b011110001100011001101101;
		13'b0001100010011: colour_data = 24'b101101011110111110110101;
		13'b0001100010100: colour_data = 24'b101101011110111110110101;
		13'b0001100010101: colour_data = 24'b101101011110111110110101;
		13'b0001100010110: colour_data = 24'b011110001100011001101101;
		13'b0001100010111: colour_data = 24'b011110001100011001101101;
		13'b0001100011000: colour_data = 24'b101101011110111110110101;
		13'b0001100011001: colour_data = 24'b101101011110111110110101;
		13'b0001100011010: colour_data = 24'b011110001100011001101101;
		13'b0001100011011: colour_data = 24'b011110001100011001101101;
		13'b0001100011100: colour_data = 24'b011110001100011001101101;
		13'b0001100011101: colour_data = 24'b101101011110111110110101;
		13'b0001100011110: colour_data = 24'b101101011110111110110101;
		13'b0001100011111: colour_data = 24'b011110001100011001101101;
		13'b0001100100000: colour_data = 24'b011110001100011001101101;
		13'b0001100100001: colour_data = 24'b101101011110111110110101;
		13'b0001100100010: colour_data = 24'b101101011110111110110101;
		13'b0001100100011: colour_data = 24'b101101011110111110110101;
		13'b0001100100100: colour_data = 24'b011110001100011001101101;
		13'b0001100100101: colour_data = 24'b011110001100011001101101;
		13'b0001100100110: colour_data = 24'b101101011110111110110101;
		13'b0001100100111: colour_data = 24'b101101011110111110110101;
		13'b0001100101000: colour_data = 24'b101101011110111110110101;
		13'b0001100101001: colour_data = 24'b011110001100011001101101;
		13'b0001100101010: colour_data = 24'b011110001100011001101101;
		13'b0001100101011: colour_data = 24'b101101011110111110110101;
		13'b0001100101100: colour_data = 24'b101101011110111110110101;
		13'b0001100101101: colour_data = 24'b011110001100011001101101;
		13'b0001100101110: colour_data = 24'b011110001100011001101101;
		13'b0001100101111: colour_data = 24'b011110001100011001101101;
		13'b0001100110000: colour_data = 24'b101101011110111110110101;
		13'b0001100110001: colour_data = 24'b101101011110111110110101;
		13'b0001100110010: colour_data = 24'b011110001100011001101101;
		13'b0001100110011: colour_data = 24'b011110001100011001101101;
		13'b0001100110100: colour_data = 24'b011010101110001101011001;
		13'b0001100110101: colour_data = 24'b101101011110111110110101;
		13'b0001100110110: colour_data = 24'b101101011110111110110101;
		13'b0001100110111: colour_data = 24'b011110001100011001101101;
		13'b0001100111000: colour_data = 24'b011110001100011001101101;
		13'b0001100111001: colour_data = 24'b101101011110111110110101;
		13'b0001100111010: colour_data = 24'b101101011110111110110101;
		13'b0001100111011: colour_data = 24'b101101011110111110110101;
		13'b0001100111100: colour_data = 24'b011110001100011001101101;
		13'b0001100111101: colour_data = 24'b011110001100011001101101;
		13'b0001100111110: colour_data = 24'b101101011110111110110101;
		13'b0001100111111: colour_data = 24'b101101011110111110110101;
		13'b0001101000000: colour_data = 24'b011110001100011001101101;
		13'b0001101000001: colour_data = 24'b011110001100011001101101;
		13'b0001101000010: colour_data = 24'b011110001100011001101101;
		13'b0001101000011: colour_data = 24'b101101011110111110110101;
		13'b0001101000100: colour_data = 24'b101101011110111110110101;
		13'b0001101000101: colour_data = 24'b011110001100011001101101;
		13'b0001101000110: colour_data = 24'b011110001100011001101101;
		13'b0001101000111: colour_data = 24'b101101011110111110110101;
		13'b0001101001000: colour_data = 24'b101101011110111110110101;
		13'b0001101001001: colour_data = 24'b101101011110111110110101;
		13'b0001101001010: colour_data = 24'b011110001100011001101101;
		13'b0001101001011: colour_data = 24'b011110001100011001101101;
		13'b0001101001100: colour_data = 24'b101101011110111110110101;
		13'b0001101001101: colour_data = 24'b101101011110111110110101;
		13'b0001101001110: colour_data = 24'b011110001100011001101101;
		13'b0001101001111: colour_data = 24'b011110001100011001101101;
		13'b0001101010000: colour_data = 24'b011110001100011001101101;
		13'b0001101010001: colour_data = 24'b101101011110111110110101;
		13'b0001101010010: colour_data = 24'b101101011110111110110101;
		13'b0001101010011: colour_data = 24'b011110001100011001101101;
		13'b0001101010100: colour_data = 24'b011110001100011001101101;
		13'b0001101010101: colour_data = 24'b011110001100011001101101;
		13'b0001101010110: colour_data = 24'b101101011110111110110101;
		13'b0001101010111: colour_data = 24'b101101011110111110110101;
		13'b0001101011000: colour_data = 24'b011110001100011001101101;
		13'b0001101011001: colour_data = 24'b011110001100011001101101;
		13'b0001101011010: colour_data = 24'b101101011110111110110101;
		13'b0001101011011: colour_data = 24'b101101011110111110110101;
		13'b0001101011100: colour_data = 24'b101101011110111110110101;
		13'b0001101011101: colour_data = 24'b011110001100011001101101;
		13'b0001101011110: colour_data = 24'b011110001100011001101101;
		13'b0001101011111: colour_data = 24'b101101011110111110110101;
		13'b0001101100000: colour_data = 24'b101101011110111110110101;
		13'b0001101100001: colour_data = 24'b011110001100011001101101;
		13'b0001101100010: colour_data = 24'b011110001100011001101101;
		13'b0001101100011: colour_data = 24'b011110001100011001101101;
		13'b0001101100100: colour_data = 24'b101101011110111110110101;
		13'b0001101100101: colour_data = 24'b101101011110111110110101;
		13'b0001101100110: colour_data = 24'b011110001100011001101101;
		13'b0001101100111: colour_data = 24'b011110001100011001101101;
		13'b0001101101000: colour_data = 24'b011110001100011001101101;
		13'b0001101101001: colour_data = 24'b101101011110111110110101;
		13'b0001101101010: colour_data = 24'b101101011110111110110101;
		13'b0001101101011: colour_data = 24'b011110001100011001101101;
		13'b0001101101100: colour_data = 24'b011110001100011001101101;
		13'b0001101101101: colour_data = 24'b101101011110111110110101;
		13'b0001101101110: colour_data = 24'b101101011110111110110101;
		13'b0001101101111: colour_data = 24'b101101011110111110110101;
		13'b0001101110000: colour_data = 24'b011110001100011001101101;
		13'b0001101110001: colour_data = 24'b011110001100011001101101;
		13'b0001101110010: colour_data = 24'b101101011110111110110101;
		13'b0001101110011: colour_data = 24'b101101011110111110110101;
		13'b0001101110100: colour_data = 24'b011110001100011001101101;
		13'b0001101110101: colour_data = 24'b011110001100011001101101;
		13'b0001101110110: colour_data = 24'b011110001100011001101101;
		13'b0001101110111: colour_data = 24'b101101011110111110110101;
		13'b0001101111000: colour_data = 24'b101101011110111110110101;
		13'b0001101111001: colour_data = 24'b011110001100011001101101;
		13'b0001101111010: colour_data = 24'b011110001100011001101101;
		13'b0001101111011: colour_data = 24'b101101011110111110110101;
		13'b0001101111100: colour_data = 24'b101101011110111110110101;
		13'b0001101111101: colour_data = 24'b101101011110111110110101;
		13'b0001101111110: colour_data = 24'b011110001100011001101101;
		13'b0001101111111: colour_data = 24'b011110001100011001101101;
		13'b0001110000000: colour_data = 24'b101101011110111110110101;
		13'b0001110000001: colour_data = 24'b101101011110111110110101;
		13'b0001110000010: colour_data = 24'b101101011110111110110101;
		13'b0001110000011: colour_data = 24'b011110001100011001101101;
		13'b0001110000100: colour_data = 24'b011110001100011001101101;
		13'b0001110000101: colour_data = 24'b101101011110111110110101;
		13'b0001110000110: colour_data = 24'b101101011110111110110101;
		13'b0001110000111: colour_data = 24'b011110001100011001101101;
		13'b0001110001000: colour_data = 24'b011110001100011001101101;
		13'b0001110001001: colour_data = 24'b001000011000111000100001;

		13'b0010000000000: colour_data = 24'b001010101100010100011000;
		13'b0010000000001: colour_data = 24'b011010101110001101011001;
		13'b0010000000010: colour_data = 24'b011010101110001101011001;
		13'b0010000000011: colour_data = 24'b001000011000111000100001;
		13'b0010000000100: colour_data = 24'b001000011000111000100001;
		13'b0010000000101: colour_data = 24'b011010101110001101011001;
		13'b0010000000110: colour_data = 24'b011010101110001101011001;
		13'b0010000000111: colour_data = 24'b001000011000111000100001;
		13'b0010000001000: colour_data = 24'b001000011000111000100001;
		13'b0010000001001: colour_data = 24'b001000011000111000100001;
		13'b0010000001010: colour_data = 24'b011010101110001101011001;
		13'b0010000001011: colour_data = 24'b011010101110001101011001;
		13'b0010000001100: colour_data = 24'b001000011000111000100001;
		13'b0010000001101: colour_data = 24'b001000011000111000100001;
		13'b0010000001110: colour_data = 24'b001000011000111000100001;
		13'b0010000001111: colour_data = 24'b011010101110001101011001;
		13'b0010000010000: colour_data = 24'b011010101110001101011001;
		13'b0010000010001: colour_data = 24'b001000011000111000100001;
		13'b0010000010010: colour_data = 24'b001000011000111000100001;
		13'b0010000010011: colour_data = 24'b011010101110001101011001;
		13'b0010000010100: colour_data = 24'b011010101110001101011001;
		13'b0010000010101: colour_data = 24'b011010101110001101011001;
		13'b0010000010110: colour_data = 24'b001000011000111000100001;
		13'b0010000010111: colour_data = 24'b001000011000111000100001;
		13'b0010000011000: colour_data = 24'b011010101110001101011001;
		13'b0010000011001: colour_data = 24'b011010101110001101011001;
		13'b0010000011010: colour_data = 24'b001000011000111000100001;
		13'b0010000011011: colour_data = 24'b001000011000111000100001;
		13'b0010000011100: colour_data = 24'b001000011000111000100001;
		13'b0010000011101: colour_data = 24'b011010101110001101011001;
		13'b0010000011110: colour_data = 24'b011010101110001101011001;
		13'b0010000011111: colour_data = 24'b001000011000111000100001;
		13'b0010000100000: colour_data = 24'b001000011000111000100001;
		13'b0010000100001: colour_data = 24'b011010101110001101011001;
		13'b0010000100010: colour_data = 24'b011010101110001101011001;
		13'b0010000100011: colour_data = 24'b011010101110001101011001;
		13'b0010000100100: colour_data = 24'b001000011000111000100001;
		13'b0010000100101: colour_data = 24'b001000011000111000100001;
		13'b0010000100110: colour_data = 24'b011010101110001101011001;
		13'b0010000100111: colour_data = 24'b011010101110001101011001;
		13'b0010000101000: colour_data = 24'b011010101110001101011001;
		13'b0010000101001: colour_data = 24'b001000011000111000100001;
		13'b0010000101010: colour_data = 24'b001000011000111000100001;
		13'b0010000101011: colour_data = 24'b011010101110001101011001;
		13'b0010000101100: colour_data = 24'b011010101110001101011001;
		13'b0010000101101: colour_data = 24'b001000011000111000100001;
		13'b0010000101110: colour_data = 24'b001000011000111000100001;
		13'b0010000101111: colour_data = 24'b001000011000111000100001;
		13'b0010000110000: colour_data = 24'b011010101110001101011001;
		13'b0010000110001: colour_data = 24'b011010101110001101011001;
		13'b0010000110010: colour_data = 24'b001000011000111000100001;
		13'b0010000110011: colour_data = 24'b001000011000111000100001;
		13'b0010000110100: colour_data = 24'b001010101100010100011000;
		13'b0010000110101: colour_data = 24'b011010101110001101011001;
		13'b0010000110110: colour_data = 24'b011010101110001101011001;
		13'b0010000110111: colour_data = 24'b001000011000111000100001;
		13'b0010000111000: colour_data = 24'b001000011000111000100001;
		13'b0010000111001: colour_data = 24'b011010101110001101011001;
		13'b0010000111010: colour_data = 24'b011010101110001101011001;
		13'b0010000111011: colour_data = 24'b011010101110001101011001;
		13'b0010000111100: colour_data = 24'b001000011000111000100001;
		13'b0010000111101: colour_data = 24'b001000011000111000100001;
		13'b0010000111110: colour_data = 24'b011010101110001101011001;
		13'b0010000111111: colour_data = 24'b011010101110001101011001;
		13'b0010001000000: colour_data = 24'b001000011000111000100001;
		13'b0010001000001: colour_data = 24'b001000011000111000100001;
		13'b0010001000010: colour_data = 24'b001000011000111000100001;
		13'b0010001000011: colour_data = 24'b011010101110001101011001;
		13'b0010001000100: colour_data = 24'b011010101110001101011001;
		13'b0010001000101: colour_data = 24'b001000011000111000100001;
		13'b0010001000110: colour_data = 24'b001000011000111000100001;
		13'b0010001000111: colour_data = 24'b011010101110001101011001;
		13'b0010001001000: colour_data = 24'b011010101110001101011001;
		13'b0010001001001: colour_data = 24'b011010101110001101011001;
		13'b0010001001010: colour_data = 24'b001000011000111000100001;
		13'b0010001001011: colour_data = 24'b001000011000111000100001;
		13'b0010001001100: colour_data = 24'b011010101110001101011001;
		13'b0010001001101: colour_data = 24'b011010101110001101011001;
		13'b0010001001110: colour_data = 24'b001000011000111000100001;
		13'b0010001001111: colour_data = 24'b001000011000111000100001;
		13'b0010001010000: colour_data = 24'b001000011000111000100001;
		13'b0010001010001: colour_data = 24'b011010101110001101011001;
		13'b0010001010010: colour_data = 24'b011010101110001101011001;
		13'b0010001010011: colour_data = 24'b001000011000111000100001;
		13'b0010001010100: colour_data = 24'b001000011000111000100001;
		13'b0010001010101: colour_data = 24'b001000011000111000100001;
		13'b0010001010110: colour_data = 24'b011010101110001101011001;
		13'b0010001010111: colour_data = 24'b011010101110001101011001;
		13'b0010001011000: colour_data = 24'b001000011000111000100001;
		13'b0010001011001: colour_data = 24'b001000011000111000100001;
		13'b0010001011010: colour_data = 24'b011010101110001101011001;
		13'b0010001011011: colour_data = 24'b011010101110001101011001;
		13'b0010001011100: colour_data = 24'b011010101110001101011001;
		13'b0010001011101: colour_data = 24'b001000011000111000100001;
		13'b0010001011110: colour_data = 24'b001000011000111000100001;
		13'b0010001011111: colour_data = 24'b011010101110001101011001;
		13'b0010001100000: colour_data = 24'b011010101110001101011001;
		13'b0010001100001: colour_data = 24'b001000011000111000100001;
		13'b0010001100010: colour_data = 24'b001000011000111000100001;
		13'b0010001100011: colour_data = 24'b001000011000111000100001;
		13'b0010001100100: colour_data = 24'b011010101110001101011001;
		13'b0010001100101: colour_data = 24'b011010101110001101011001;
		13'b0010001100110: colour_data = 24'b001000011000111000100001;
		13'b0010001100111: colour_data = 24'b001000011000111000100001;
		13'b0010001101000: colour_data = 24'b001000011000111000100001;
		13'b0010001101001: colour_data = 24'b011010101110001101011001;
		13'b0010001101010: colour_data = 24'b011010101110001101011001;
		13'b0010001101011: colour_data = 24'b001000011000111000100001;
		13'b0010001101100: colour_data = 24'b001000011000111000100001;
		13'b0010001101101: colour_data = 24'b011010101110001101011001;
		13'b0010001101110: colour_data = 24'b011010101110001101011001;
		13'b0010001101111: colour_data = 24'b011010101110001101011001;
		13'b0010001110000: colour_data = 24'b001000011000111000100001;
		13'b0010001110001: colour_data = 24'b001000011000111000100001;
		13'b0010001110010: colour_data = 24'b011010101110001101011001;
		13'b0010001110011: colour_data = 24'b011010101110001101011001;
		13'b0010001110100: colour_data = 24'b001000011000111000100001;
		13'b0010001110101: colour_data = 24'b001000011000111000100001;
		13'b0010001110110: colour_data = 24'b001000011000111000100001;
		13'b0010001110111: colour_data = 24'b011010101110001101011001;
		13'b0010001111000: colour_data = 24'b011010101110001101011001;
		13'b0010001111001: colour_data = 24'b001000011000111000100001;
		13'b0010001111010: colour_data = 24'b001000011000111000100001;
		13'b0010001111011: colour_data = 24'b011010101110001101011001;
		13'b0010001111100: colour_data = 24'b011010101110001101011001;
		13'b0010001111101: colour_data = 24'b011010101110001101011001;
		13'b0010001111110: colour_data = 24'b001000011000111000100001;
		13'b0010001111111: colour_data = 24'b001000011000111000100001;
		13'b0010010000000: colour_data = 24'b011010101110001101011001;
		13'b0010010000001: colour_data = 24'b011010101110001101011001;
		13'b0010010000010: colour_data = 24'b011010101110001101011001;
		13'b0010010000011: colour_data = 24'b001000011000111000100001;
		13'b0010010000100: colour_data = 24'b001000011000111000100001;
		13'b0010010000101: colour_data = 24'b011010101110001101011001;
		13'b0010010000110: colour_data = 24'b011010101110001101011001;
		13'b0010010000111: colour_data = 24'b001000011000111000100001;
		13'b0010010001000: colour_data = 24'b001000011000111000100001;
		13'b0010010001001: colour_data = 24'b000110000110110100011000;

		13'b0010100000000: colour_data = 24'b001010101100010100011000;
		13'b0010100000001: colour_data = 24'b011010101110001101011001;
		13'b0010100000010: colour_data = 24'b011010101110001101011001;
		13'b0010100000011: colour_data = 24'b001000011000111000100001;
		13'b0010100000100: colour_data = 24'b001000011000111000100001;
		13'b0010100000101: colour_data = 24'b011010101110001101011001;
		13'b0010100000110: colour_data = 24'b011010101110001101011001;
		13'b0010100000111: colour_data = 24'b001000011000111000100001;
		13'b0010100001000: colour_data = 24'b001000011000111000100001;
		13'b0010100001001: colour_data = 24'b001000011000111000100001;
		13'b0010100001010: colour_data = 24'b011010101110001101011001;
		13'b0010100001011: colour_data = 24'b011010101110001101011001;
		13'b0010100001100: colour_data = 24'b001000011000111000100001;
		13'b0010100001101: colour_data = 24'b001000011000111000100001;
		13'b0010100001110: colour_data = 24'b001000011000111000100001;
		13'b0010100001111: colour_data = 24'b011010101110001101011001;
		13'b0010100010000: colour_data = 24'b011010101110001101011001;
		13'b0010100010001: colour_data = 24'b001000011000111000100001;
		13'b0010100010010: colour_data = 24'b001000011000111000100001;
		13'b0010100010011: colour_data = 24'b011010101110001101011001;
		13'b0010100010100: colour_data = 24'b011010101110001101011001;
		13'b0010100010101: colour_data = 24'b011010101110001101011001;
		13'b0010100010110: colour_data = 24'b001000011000111000100001;
		13'b0010100010111: colour_data = 24'b001000011000111000100001;
		13'b0010100011000: colour_data = 24'b011010101110001101011001;
		13'b0010100011001: colour_data = 24'b011010101110001101011001;
		13'b0010100011010: colour_data = 24'b001000011000111000100001;
		13'b0010100011011: colour_data = 24'b001000011000111000100001;
		13'b0010100011100: colour_data = 24'b001000011000111000100001;
		13'b0010100011101: colour_data = 24'b011010101110001101011001;
		13'b0010100011110: colour_data = 24'b011010101110001101011001;
		13'b0010100011111: colour_data = 24'b001000011000111000100001;
		13'b0010100100000: colour_data = 24'b001000011000111000100001;
		13'b0010100100001: colour_data = 24'b011010101110001101011001;
		13'b0010100100010: colour_data = 24'b011010101110001101011001;
		13'b0010100100011: colour_data = 24'b011010101110001101011001;
		13'b0010100100100: colour_data = 24'b001000011000111000100001;
		13'b0010100100101: colour_data = 24'b001000011000111000100001;
		13'b0010100100110: colour_data = 24'b011010101110001101011001;
		13'b0010100100111: colour_data = 24'b011010101110001101011001;
		13'b0010100101000: colour_data = 24'b011010101110001101011001;
		13'b0010100101001: colour_data = 24'b001000011000111000100001;
		13'b0010100101010: colour_data = 24'b001000011000111000100001;
		13'b0010100101011: colour_data = 24'b011010101110001101011001;
		13'b0010100101100: colour_data = 24'b011010101110001101011001;
		13'b0010100101101: colour_data = 24'b001000011000111000100001;
		13'b0010100101110: colour_data = 24'b001000011000111000100001;
		13'b0010100101111: colour_data = 24'b001000011000111000100001;
		13'b0010100110000: colour_data = 24'b011010101110001101011001;
		13'b0010100110001: colour_data = 24'b011010101110001101011001;
		13'b0010100110010: colour_data = 24'b001000011000111000100001;
		13'b0010100110011: colour_data = 24'b001000011000111000100001;
		13'b0010100110100: colour_data = 24'b001010101100010100011000;
		13'b0010100110101: colour_data = 24'b011010101110001101011001;
		13'b0010100110110: colour_data = 24'b011010101110001101011001;
		13'b0010100110111: colour_data = 24'b001000011000111000100001;
		13'b0010100111000: colour_data = 24'b001000011000111000100001;
		13'b0010100111001: colour_data = 24'b011010101110001101011001;
		13'b0010100111010: colour_data = 24'b011010101110001101011001;
		13'b0010100111011: colour_data = 24'b011010101110001101011001;
		13'b0010100111100: colour_data = 24'b001000011000111000100001;
		13'b0010100111101: colour_data = 24'b001000011000111000100001;
		13'b0010100111110: colour_data = 24'b011010101110001101011001;
		13'b0010100111111: colour_data = 24'b011010101110001101011001;
		13'b0010101000000: colour_data = 24'b001000011000111000100001;
		13'b0010101000001: colour_data = 24'b001000011000111000100001;
		13'b0010101000010: colour_data = 24'b001000011000111000100001;
		13'b0010101000011: colour_data = 24'b011010101110001101011001;
		13'b0010101000100: colour_data = 24'b011010101110001101011001;
		13'b0010101000101: colour_data = 24'b001000011000111000100001;
		13'b0010101000110: colour_data = 24'b001000011000111000100001;
		13'b0010101000111: colour_data = 24'b011010101110001101011001;
		13'b0010101001000: colour_data = 24'b011010101110001101011001;
		13'b0010101001001: colour_data = 24'b011010101110001101011001;
		13'b0010101001010: colour_data = 24'b001000011000111000100001;
		13'b0010101001011: colour_data = 24'b001000011000111000100001;
		13'b0010101001100: colour_data = 24'b011010101110001101011001;
		13'b0010101001101: colour_data = 24'b011010101110001101011001;
		13'b0010101001110: colour_data = 24'b001000011000111000100001;
		13'b0010101001111: colour_data = 24'b001000011000111000100001;
		13'b0010101010000: colour_data = 24'b001000011000111000100001;
		13'b0010101010001: colour_data = 24'b011010101110001101011001;
		13'b0010101010010: colour_data = 24'b011010101110001101011001;
		13'b0010101010011: colour_data = 24'b001000011000111000100001;
		13'b0010101010100: colour_data = 24'b001000011000111000100001;
		13'b0010101010101: colour_data = 24'b001000011000111000100001;
		13'b0010101010110: colour_data = 24'b011010101110001101011001;
		13'b0010101010111: colour_data = 24'b011010101110001101011001;
		13'b0010101011000: colour_data = 24'b001000011000111000100001;
		13'b0010101011001: colour_data = 24'b001000011000111000100001;
		13'b0010101011010: colour_data = 24'b011010101110001101011001;
		13'b0010101011011: colour_data = 24'b011010101110001101011001;
		13'b0010101011100: colour_data = 24'b011010101110001101011001;
		13'b0010101011101: colour_data = 24'b001000011000111000100001;
		13'b0010101011110: colour_data = 24'b001000011000111000100001;
		13'b0010101011111: colour_data = 24'b011010101110001101011001;
		13'b0010101100000: colour_data = 24'b011010101110001101011001;
		13'b0010101100001: colour_data = 24'b001000011000111000100001;
		13'b0010101100010: colour_data = 24'b001000011000111000100001;
		13'b0010101100011: colour_data = 24'b001000011000111000100001;
		13'b0010101100100: colour_data = 24'b011010101110001101011001;
		13'b0010101100101: colour_data = 24'b011010101110001101011001;
		13'b0010101100110: colour_data = 24'b001000011000111000100001;
		13'b0010101100111: colour_data = 24'b001000011000111000100001;
		13'b0010101101000: colour_data = 24'b001000011000111000100001;
		13'b0010101101001: colour_data = 24'b011010101110001101011001;
		13'b0010101101010: colour_data = 24'b011010101110001101011001;
		13'b0010101101011: colour_data = 24'b001000011000111000100001;
		13'b0010101101100: colour_data = 24'b001000011000111000100001;
		13'b0010101101101: colour_data = 24'b011010101110001101011001;
		13'b0010101101110: colour_data = 24'b011010101110001101011001;
		13'b0010101101111: colour_data = 24'b011010101110001101011001;
		13'b0010101110000: colour_data = 24'b001000011000111000100001;
		13'b0010101110001: colour_data = 24'b001000011000111000100001;
		13'b0010101110010: colour_data = 24'b011010101110001101011001;
		13'b0010101110011: colour_data = 24'b011010101110001101011001;
		13'b0010101110100: colour_data = 24'b001000011000111000100001;
		13'b0010101110101: colour_data = 24'b001000011000111000100001;
		13'b0010101110110: colour_data = 24'b001000011000111000100001;
		13'b0010101110111: colour_data = 24'b011010101110001101011001;
		13'b0010101111000: colour_data = 24'b011010101110001101011001;
		13'b0010101111001: colour_data = 24'b001000011000111000100001;
		13'b0010101111010: colour_data = 24'b001000011000111000100001;
		13'b0010101111011: colour_data = 24'b011010101110001101011001;
		13'b0010101111100: colour_data = 24'b011010101110001101011001;
		13'b0010101111101: colour_data = 24'b011010101110001101011001;
		13'b0010101111110: colour_data = 24'b001000011000111000100001;
		13'b0010101111111: colour_data = 24'b001000011000111000100001;
		13'b0010110000000: colour_data = 24'b011010101110001101011001;
		13'b0010110000001: colour_data = 24'b011010101110001101011001;
		13'b0010110000010: colour_data = 24'b011010101110001101011001;
		13'b0010110000011: colour_data = 24'b001000011000111000100001;
		13'b0010110000100: colour_data = 24'b001000011000111000100001;
		13'b0010110000101: colour_data = 24'b011010101110001101011001;
		13'b0010110000110: colour_data = 24'b011010101110001101011001;
		13'b0010110000111: colour_data = 24'b001000011000111000100001;
		13'b0010110001000: colour_data = 24'b001000011000111000100001;
		13'b0010110001001: colour_data = 24'b000110000110110100011000;

		13'b0011000000000: colour_data = 24'b001010101100010100011000;
		13'b0011000000001: colour_data = 24'b011010101110001101011001;
		13'b0011000000010: colour_data = 24'b011010101110001101011001;
		13'b0011000000011: colour_data = 24'b001000011000111000100001;
		13'b0011000000100: colour_data = 24'b001000011000111000100001;
		13'b0011000000101: colour_data = 24'b011010101110001101011001;
		13'b0011000000110: colour_data = 24'b011010101110001101011001;
		13'b0011000000111: colour_data = 24'b001000011000111000100001;
		13'b0011000001000: colour_data = 24'b001000011000111000100001;
		13'b0011000001001: colour_data = 24'b001000011000111000100001;
		13'b0011000001010: colour_data = 24'b011010101110001101011001;
		13'b0011000001011: colour_data = 24'b011010101110001101011001;
		13'b0011000001100: colour_data = 24'b001000011000111000100001;
		13'b0011000001101: colour_data = 24'b000110000110110100011000;
		13'b0011000001110: colour_data = 24'b001000011000111000100001;
		13'b0011000001111: colour_data = 24'b011010101110001101011001;
		13'b0011000010000: colour_data = 24'b011010101110001101011001;
		13'b0011000010001: colour_data = 24'b001000011000111000100001;
		13'b0011000010010: colour_data = 24'b000110000110110100011000;
		13'b0011000010011: colour_data = 24'b011010101110001101011001;
		13'b0011000010100: colour_data = 24'b011010101110001101011001;
		13'b0011000010101: colour_data = 24'b011010101110001101011001;
		13'b0011000010110: colour_data = 24'b001000011000111000100001;
		13'b0011000010111: colour_data = 24'b001000011000111000100001;
		13'b0011000011000: colour_data = 24'b011010101110001101011001;
		13'b0011000011001: colour_data = 24'b011010101110001101011001;
		13'b0011000011010: colour_data = 24'b001000011000111000100001;
		13'b0011000011011: colour_data = 24'b001000011000111000100001;
		13'b0011000011100: colour_data = 24'b001000011000111000100001;
		13'b0011000011101: colour_data = 24'b011010101110001101011001;
		13'b0011000011110: colour_data = 24'b011010101110001101011001;
		13'b0011000011111: colour_data = 24'b001000011000111000100001;
		13'b0011000100000: colour_data = 24'b000110000110110100011000;
		13'b0011000100001: colour_data = 24'b011010101110001101011001;
		13'b0011000100010: colour_data = 24'b011010101110001101011001;
		13'b0011000100011: colour_data = 24'b011010101110001101011001;
		13'b0011000100100: colour_data = 24'b001000011000111000100001;
		13'b0011000100101: colour_data = 24'b000110000110110100011000;
		13'b0011000100110: colour_data = 24'b011010101110001101011001;
		13'b0011000100111: colour_data = 24'b011010101110001101011001;
		13'b0011000101000: colour_data = 24'b011010101110001101011001;
		13'b0011000101001: colour_data = 24'b001000011000111000100001;
		13'b0011000101010: colour_data = 24'b001000011000111000100001;
		13'b0011000101011: colour_data = 24'b011010101110001101011001;
		13'b0011000101100: colour_data = 24'b011010101110001101011001;
		13'b0011000101101: colour_data = 24'b001000011000111000100001;
		13'b0011000101110: colour_data = 24'b001000011000111000100001;
		13'b0011000101111: colour_data = 24'b001000011000111000100001;
		13'b0011000110000: colour_data = 24'b011010101110001101011001;
		13'b0011000110001: colour_data = 24'b011010101110001101011001;
		13'b0011000110010: colour_data = 24'b001000011000111000100001;
		13'b0011000110011: colour_data = 24'b000110000110110100011000;
		13'b0011000110100: colour_data = 24'b001010101100010100011000;
		13'b0011000110101: colour_data = 24'b011010101110001101011001;
		13'b0011000110110: colour_data = 24'b011010101110001101011001;
		13'b0011000110111: colour_data = 24'b001000011000111000100001;
		13'b0011000111000: colour_data = 24'b000110000110110100011000;
		13'b0011000111001: colour_data = 24'b011010101110001101011001;
		13'b0011000111010: colour_data = 24'b011010101110001101011001;
		13'b0011000111011: colour_data = 24'b011010101110001101011001;
		13'b0011000111100: colour_data = 24'b001000011000111000100001;
		13'b0011000111101: colour_data = 24'b001000011000111000100001;
		13'b0011000111110: colour_data = 24'b011010101110001101011001;
		13'b0011000111111: colour_data = 24'b011010101110001101011001;
		13'b0011001000000: colour_data = 24'b001000011000111000100001;
		13'b0011001000001: colour_data = 24'b000110000110110100011000;
		13'b0011001000010: colour_data = 24'b001000011000111000100001;
		13'b0011001000011: colour_data = 24'b011010101110001101011001;
		13'b0011001000100: colour_data = 24'b011010101110001101011001;
		13'b0011001000101: colour_data = 24'b001000011000111000100001;
		13'b0011001000110: colour_data = 24'b000110000110110100011000;
		13'b0011001000111: colour_data = 24'b011010101110001101011001;
		13'b0011001001000: colour_data = 24'b011010101110001101011001;
		13'b0011001001001: colour_data = 24'b011010101110001101011001;
		13'b0011001001010: colour_data = 24'b001000011000111000100001;
		13'b0011001001011: colour_data = 24'b000110000110110100011000;
		13'b0011001001100: colour_data = 24'b011010101110001101011001;
		13'b0011001001101: colour_data = 24'b011010101110001101011001;
		13'b0011001001110: colour_data = 24'b001000011000111000100001;
		13'b0011001001111: colour_data = 24'b001000011000111000100001;
		13'b0011001010000: colour_data = 24'b001000011000111000100001;
		13'b0011001010001: colour_data = 24'b011010101110001101011001;
		13'b0011001010010: colour_data = 24'b011010101110001101011001;
		13'b0011001010011: colour_data = 24'b001000011000111000100001;
		13'b0011001010100: colour_data = 24'b000110000110110100011000;
		13'b0011001010101: colour_data = 24'b001000011000111000100001;
		13'b0011001010110: colour_data = 24'b011010101110001101011001;
		13'b0011001010111: colour_data = 24'b011010101110001101011001;
		13'b0011001011000: colour_data = 24'b001000011000111000100001;
		13'b0011001011001: colour_data = 24'b000110000110110100011000;
		13'b0011001011010: colour_data = 24'b011010101110001101011001;
		13'b0011001011011: colour_data = 24'b011010101110001101011001;
		13'b0011001011100: colour_data = 24'b011010101110001101011001;
		13'b0011001011101: colour_data = 24'b001000011000111000100001;
		13'b0011001011110: colour_data = 24'b001000011000111000100001;
		13'b0011001011111: colour_data = 24'b011010101110001101011001;
		13'b0011001100000: colour_data = 24'b011010101110001101011001;
		13'b0011001100001: colour_data = 24'b001000011000111000100001;
		13'b0011001100010: colour_data = 24'b001000011000111000100001;
		13'b0011001100011: colour_data = 24'b001000011000111000100001;
		13'b0011001100100: colour_data = 24'b011010101110001101011001;
		13'b0011001100101: colour_data = 24'b011010101110001101011001;
		13'b0011001100110: colour_data = 24'b001000011000111000100001;
		13'b0011001100111: colour_data = 24'b000110000110110100011000;
		13'b0011001101000: colour_data = 24'b001000011000111000100001;
		13'b0011001101001: colour_data = 24'b011010101110001101011001;
		13'b0011001101010: colour_data = 24'b011010101110001101011001;
		13'b0011001101011: colour_data = 24'b001000011000111000100001;
		13'b0011001101100: colour_data = 24'b000110000110110100011000;
		13'b0011001101101: colour_data = 24'b011010101110001101011001;
		13'b0011001101110: colour_data = 24'b011010101110001101011001;
		13'b0011001101111: colour_data = 24'b011010101110001101011001;
		13'b0011001110000: colour_data = 24'b001000011000111000100001;
		13'b0011001110001: colour_data = 24'b001000011000111000100001;
		13'b0011001110010: colour_data = 24'b011010101110001101011001;
		13'b0011001110011: colour_data = 24'b011010101110001101011001;
		13'b0011001110100: colour_data = 24'b001000011000111000100001;
		13'b0011001110101: colour_data = 24'b001000011000111000100001;
		13'b0011001110110: colour_data = 24'b001000011000111000100001;
		13'b0011001110111: colour_data = 24'b011010101110001101011001;
		13'b0011001111000: colour_data = 24'b011010101110001101011001;
		13'b0011001111001: colour_data = 24'b001000011000111000100001;
		13'b0011001111010: colour_data = 24'b000110000110110100011000;
		13'b0011001111011: colour_data = 24'b011010101110001101011001;
		13'b0011001111100: colour_data = 24'b011010101110001101011001;
		13'b0011001111101: colour_data = 24'b011010101110001101011001;
		13'b0011001111110: colour_data = 24'b001000011000111000100001;
		13'b0011001111111: colour_data = 24'b000110000110110100011000;
		13'b0011010000000: colour_data = 24'b011010101110001101011001;
		13'b0011010000001: colour_data = 24'b011010101110001101011001;
		13'b0011010000010: colour_data = 24'b011010101110001101011001;
		13'b0011010000011: colour_data = 24'b001000011000111000100001;
		13'b0011010000100: colour_data = 24'b001000011000111000100001;
		13'b0011010000101: colour_data = 24'b011010101110001101011001;
		13'b0011010000110: colour_data = 24'b011010101110001101011001;
		13'b0011010000111: colour_data = 24'b001000011000111000100001;
		13'b0011010001000: colour_data = 24'b000110000110110100011000;
		13'b0011010001001: colour_data = 24'b000110000110110100011000;

		13'b0011100000000: colour_data = 24'b001010101100010100011000;
		13'b0011100000001: colour_data = 24'b011010101110001101011001;
		13'b0011100000010: colour_data = 24'b011010101110001101011001;
		13'b0011100000011: colour_data = 24'b001000011000111000100001;
		13'b0011100000100: colour_data = 24'b001000011000111000100001;
		13'b0011100000101: colour_data = 24'b011010101110001101011001;
		13'b0011100000110: colour_data = 24'b011010101110001101011001;
		13'b0011100000111: colour_data = 24'b001000011000111000100001;
		13'b0011100001000: colour_data = 24'b001000011000111000100001;
		13'b0011100001001: colour_data = 24'b001000011000111000100001;
		13'b0011100001010: colour_data = 24'b011010101110001101011001;
		13'b0011100001011: colour_data = 24'b011010101110001101011001;
		13'b0011100001100: colour_data = 24'b001000011000111000100001;
		13'b0011100001101: colour_data = 24'b000110000110110100011000;
		13'b0011100001110: colour_data = 24'b001000011000111000100001;
		13'b0011100001111: colour_data = 24'b011010101110001101011001;
		13'b0011100010000: colour_data = 24'b011010101110001101011001;
		13'b0011100010001: colour_data = 24'b001000011000111000100001;
		13'b0011100010010: colour_data = 24'b000110000110110100011000;
		13'b0011100010011: colour_data = 24'b011010101110001101011001;
		13'b0011100010100: colour_data = 24'b011010101110001101011001;
		13'b0011100010101: colour_data = 24'b011010101110001101011001;
		13'b0011100010110: colour_data = 24'b001000011000111000100001;
		13'b0011100010111: colour_data = 24'b001000011000111000100001;
		13'b0011100011000: colour_data = 24'b011010101110001101011001;
		13'b0011100011001: colour_data = 24'b011010101110001101011001;
		13'b0011100011010: colour_data = 24'b001000011000111000100001;
		13'b0011100011011: colour_data = 24'b001000011000111000100001;
		13'b0011100011100: colour_data = 24'b001000011000111000100001;
		13'b0011100011101: colour_data = 24'b011010101110001101011001;
		13'b0011100011110: colour_data = 24'b011010101110001101011001;
		13'b0011100011111: colour_data = 24'b001000011000111000100001;
		13'b0011100100000: colour_data = 24'b000110000110110100011000;
		13'b0011100100001: colour_data = 24'b011010101110001101011001;
		13'b0011100100010: colour_data = 24'b011010101110001101011001;
		13'b0011100100011: colour_data = 24'b011010101110001101011001;
		13'b0011100100100: colour_data = 24'b001000011000111000100001;
		13'b0011100100101: colour_data = 24'b000110000110110100011000;
		13'b0011100100110: colour_data = 24'b011010101110001101011001;
		13'b0011100100111: colour_data = 24'b011010101110001101011001;
		13'b0011100101000: colour_data = 24'b011010101110001101011001;
		13'b0011100101001: colour_data = 24'b001000011000111000100001;
		13'b0011100101010: colour_data = 24'b001000011000111000100001;
		13'b0011100101011: colour_data = 24'b011010101110001101011001;
		13'b0011100101100: colour_data = 24'b011010101110001101011001;
		13'b0011100101101: colour_data = 24'b001000011000111000100001;
		13'b0011100101110: colour_data = 24'b001000011000111000100001;
		13'b0011100101111: colour_data = 24'b001000011000111000100001;
		13'b0011100110000: colour_data = 24'b011010101110001101011001;
		13'b0011100110001: colour_data = 24'b011010101110001101011001;
		13'b0011100110010: colour_data = 24'b001000011000111000100001;
		13'b0011100110011: colour_data = 24'b000110000110110100011000;
		13'b0011100110100: colour_data = 24'b001010101100010100011000;
		13'b0011100110101: colour_data = 24'b011010101110001101011001;
		13'b0011100110110: colour_data = 24'b011010101110001101011001;
		13'b0011100110111: colour_data = 24'b001000011000111000100001;
		13'b0011100111000: colour_data = 24'b000110000110110100011000;
		13'b0011100111001: colour_data = 24'b011010101110001101011001;
		13'b0011100111010: colour_data = 24'b011010101110001101011001;
		13'b0011100111011: colour_data = 24'b011010101110001101011001;
		13'b0011100111100: colour_data = 24'b001000011000111000100001;
		13'b0011100111101: colour_data = 24'b001000011000111000100001;
		13'b0011100111110: colour_data = 24'b011010101110001101011001;
		13'b0011100111111: colour_data = 24'b011010101110001101011001;
		13'b0011101000000: colour_data = 24'b001000011000111000100001;
		13'b0011101000001: colour_data = 24'b000110000110110100011000;
		13'b0011101000010: colour_data = 24'b001000011000111000100001;
		13'b0011101000011: colour_data = 24'b011010101110001101011001;
		13'b0011101000100: colour_data = 24'b011010101110001101011001;
		13'b0011101000101: colour_data = 24'b001000011000111000100001;
		13'b0011101000110: colour_data = 24'b000110000110110100011000;
		13'b0011101000111: colour_data = 24'b011010101110001101011001;
		13'b0011101001000: colour_data = 24'b011010101110001101011001;
		13'b0011101001001: colour_data = 24'b011010101110001101011001;
		13'b0011101001010: colour_data = 24'b001000011000111000100001;
		13'b0011101001011: colour_data = 24'b000110000110110100011000;
		13'b0011101001100: colour_data = 24'b011010101110001101011001;
		13'b0011101001101: colour_data = 24'b011010101110001101011001;
		13'b0011101001110: colour_data = 24'b001000011000111000100001;
		13'b0011101001111: colour_data = 24'b001000011000111000100001;
		13'b0011101010000: colour_data = 24'b001000011000111000100001;
		13'b0011101010001: colour_data = 24'b011010101110001101011001;
		13'b0011101010010: colour_data = 24'b011010101110001101011001;
		13'b0011101010011: colour_data = 24'b001000011000111000100001;
		13'b0011101010100: colour_data = 24'b000110000110110100011000;
		13'b0011101010101: colour_data = 24'b001000011000111000100001;
		13'b0011101010110: colour_data = 24'b011010101110001101011001;
		13'b0011101010111: colour_data = 24'b011010101110001101011001;
		13'b0011101011000: colour_data = 24'b001000011000111000100001;
		13'b0011101011001: colour_data = 24'b000110000110110100011000;
		13'b0011101011010: colour_data = 24'b011010101110001101011001;
		13'b0011101011011: colour_data = 24'b011010101110001101011001;
		13'b0011101011100: colour_data = 24'b011010101110001101011001;
		13'b0011101011101: colour_data = 24'b001000011000111000100001;
		13'b0011101011110: colour_data = 24'b001000011000111000100001;
		13'b0011101011111: colour_data = 24'b011010101110001101011001;
		13'b0011101100000: colour_data = 24'b011010101110001101011001;
		13'b0011101100001: colour_data = 24'b001000011000111000100001;
		13'b0011101100010: colour_data = 24'b001000011000111000100001;
		13'b0011101100011: colour_data = 24'b001000011000111000100001;
		13'b0011101100100: colour_data = 24'b011010101110001101011001;
		13'b0011101100101: colour_data = 24'b011010101110001101011001;
		13'b0011101100110: colour_data = 24'b001000011000111000100001;
		13'b0011101100111: colour_data = 24'b000110000110110100011000;
		13'b0011101101000: colour_data = 24'b001000011000111000100001;
		13'b0011101101001: colour_data = 24'b011010101110001101011001;
		13'b0011101101010: colour_data = 24'b011010101110001101011001;
		13'b0011101101011: colour_data = 24'b001000011000111000100001;
		13'b0011101101100: colour_data = 24'b000110000110110100011000;
		13'b0011101101101: colour_data = 24'b011010101110001101011001;
		13'b0011101101110: colour_data = 24'b011010101110001101011001;
		13'b0011101101111: colour_data = 24'b011010101110001101011001;
		13'b0011101110000: colour_data = 24'b001000011000111000100001;
		13'b0011101110001: colour_data = 24'b001000011000111000100001;
		13'b0011101110010: colour_data = 24'b011010101110001101011001;
		13'b0011101110011: colour_data = 24'b011010101110001101011001;
		13'b0011101110100: colour_data = 24'b001000011000111000100001;
		13'b0011101110101: colour_data = 24'b001000011000111000100001;
		13'b0011101110110: colour_data = 24'b001000011000111000100001;
		13'b0011101110111: colour_data = 24'b011010101110001101011001;
		13'b0011101111000: colour_data = 24'b011010101110001101011001;
		13'b0011101111001: colour_data = 24'b001000011000111000100001;
		13'b0011101111010: colour_data = 24'b000110000110110100011000;
		13'b0011101111011: colour_data = 24'b011010101110001101011001;
		13'b0011101111100: colour_data = 24'b011010101110001101011001;
		13'b0011101111101: colour_data = 24'b011010101110001101011001;
		13'b0011101111110: colour_data = 24'b001000011000111000100001;
		13'b0011101111111: colour_data = 24'b000110000110110100011000;
		13'b0011110000000: colour_data = 24'b011010101110001101011001;
		13'b0011110000001: colour_data = 24'b011010101110001101011001;
		13'b0011110000010: colour_data = 24'b011010101110001101011001;
		13'b0011110000011: colour_data = 24'b001000011000111000100001;
		13'b0011110000100: colour_data = 24'b001000011000111000100001;
		13'b0011110000101: colour_data = 24'b011010101110001101011001;
		13'b0011110000110: colour_data = 24'b011010101110001101011001;
		13'b0011110000111: colour_data = 24'b001000011000111000100001;
		13'b0011110001000: colour_data = 24'b000110000110110100011000;
		13'b0011110001001: colour_data = 24'b000110000110110100011000;

		13'b0100000000000: colour_data = 24'b001010101100010100011000;
		13'b0100000000001: colour_data = 24'b011010101110001101011001;
		13'b0100000000010: colour_data = 24'b011010101110001101011001;
		13'b0100000000011: colour_data = 24'b001000011000111000100001;
		13'b0100000000100: colour_data = 24'b001000011000111000100001;
		13'b0100000000101: colour_data = 24'b011010101110001101011001;
		13'b0100000000110: colour_data = 24'b011010101110001101011001;
		13'b0100000000111: colour_data = 24'b001000011000111000100001;
		13'b0100000001000: colour_data = 24'b001000011000111000100001;
		13'b0100000001001: colour_data = 24'b001000011000111000100001;
		13'b0100000001010: colour_data = 24'b011010101110001101011001;
		13'b0100000001011: colour_data = 24'b011010101110001101011001;
		13'b0100000001100: colour_data = 24'b001000011000111000100001;
		13'b0100000001101: colour_data = 24'b000110000110110100011000;
		13'b0100000001110: colour_data = 24'b001000011000111000100001;
		13'b0100000001111: colour_data = 24'b011010101110001101011001;
		13'b0100000010000: colour_data = 24'b011010101110001101011001;
		13'b0100000010001: colour_data = 24'b001000011000111000100001;
		13'b0100000010010: colour_data = 24'b000110000110110100011000;
		13'b0100000010011: colour_data = 24'b011010101110001101011001;
		13'b0100000010100: colour_data = 24'b011010101110001101011001;
		13'b0100000010101: colour_data = 24'b011010101110001101011001;
		13'b0100000010110: colour_data = 24'b001000011000111000100001;
		13'b0100000010111: colour_data = 24'b001000011000111000100001;
		13'b0100000011000: colour_data = 24'b011010101110001101011001;
		13'b0100000011001: colour_data = 24'b011010101110001101011001;
		13'b0100000011010: colour_data = 24'b001000011000111000100001;
		13'b0100000011011: colour_data = 24'b001000011000111000100001;
		13'b0100000011100: colour_data = 24'b001000011000111000100001;
		13'b0100000011101: colour_data = 24'b011010101110001101011001;
		13'b0100000011110: colour_data = 24'b011010101110001101011001;
		13'b0100000011111: colour_data = 24'b001000011000111000100001;
		13'b0100000100000: colour_data = 24'b000110000110110100011000;
		13'b0100000100001: colour_data = 24'b011010101110001101011001;
		13'b0100000100010: colour_data = 24'b011010101110001101011001;
		13'b0100000100011: colour_data = 24'b011010101110001101011001;
		13'b0100000100100: colour_data = 24'b001000011000111000100001;
		13'b0100000100101: colour_data = 24'b000110000110110100011000;
		13'b0100000100110: colour_data = 24'b011010101110001101011001;
		13'b0100000100111: colour_data = 24'b011010101110001101011001;
		13'b0100000101000: colour_data = 24'b011010101110001101011001;
		13'b0100000101001: colour_data = 24'b001000011000111000100001;
		13'b0100000101010: colour_data = 24'b001000011000111000100001;
		13'b0100000101011: colour_data = 24'b011010101110001101011001;
		13'b0100000101100: colour_data = 24'b011010101110001101011001;
		13'b0100000101101: colour_data = 24'b001000011000111000100001;
		13'b0100000101110: colour_data = 24'b001000011000111000100001;
		13'b0100000101111: colour_data = 24'b001000011000111000100001;
		13'b0100000110000: colour_data = 24'b011010101110001101011001;
		13'b0100000110001: colour_data = 24'b011010101110001101011001;
		13'b0100000110010: colour_data = 24'b001000011000111000100001;
		13'b0100000110011: colour_data = 24'b000110000110110100011000;
		13'b0100000110100: colour_data = 24'b001010101100010100011000;
		13'b0100000110101: colour_data = 24'b011010101110001101011001;
		13'b0100000110110: colour_data = 24'b011010101110001101011001;
		13'b0100000110111: colour_data = 24'b001000011000111000100001;
		13'b0100000111000: colour_data = 24'b000110000110110100011000;
		13'b0100000111001: colour_data = 24'b011010101110001101011001;
		13'b0100000111010: colour_data = 24'b011010101110001101011001;
		13'b0100000111011: colour_data = 24'b011010101110001101011001;
		13'b0100000111100: colour_data = 24'b001000011000111000100001;
		13'b0100000111101: colour_data = 24'b001000011000111000100001;
		13'b0100000111110: colour_data = 24'b011010101110001101011001;
		13'b0100000111111: colour_data = 24'b011010101110001101011001;
		13'b0100001000000: colour_data = 24'b001000011000111000100001;
		13'b0100001000001: colour_data = 24'b000110000110110100011000;
		13'b0100001000010: colour_data = 24'b001000011000111000100001;
		13'b0100001000011: colour_data = 24'b011010101110001101011001;
		13'b0100001000100: colour_data = 24'b011010101110001101011001;
		13'b0100001000101: colour_data = 24'b001000011000111000100001;
		13'b0100001000110: colour_data = 24'b000110000110110100011000;
		13'b0100001000111: colour_data = 24'b011010101110001101011001;
		13'b0100001001000: colour_data = 24'b011010101110001101011001;
		13'b0100001001001: colour_data = 24'b011010101110001101011001;
		13'b0100001001010: colour_data = 24'b001000011000111000100001;
		13'b0100001001011: colour_data = 24'b000110000110110100011000;
		13'b0100001001100: colour_data = 24'b011010101110001101011001;
		13'b0100001001101: colour_data = 24'b011010101110001101011001;
		13'b0100001001110: colour_data = 24'b001000011000111000100001;
		13'b0100001001111: colour_data = 24'b001000011000111000100001;
		13'b0100001010000: colour_data = 24'b001000011000111000100001;
		13'b0100001010001: colour_data = 24'b011010101110001101011001;
		13'b0100001010010: colour_data = 24'b011010101110001101011001;
		13'b0100001010011: colour_data = 24'b001000011000111000100001;
		13'b0100001010100: colour_data = 24'b000110000110110100011000;
		13'b0100001010101: colour_data = 24'b001000011000111000100001;
		13'b0100001010110: colour_data = 24'b011010101110001101011001;
		13'b0100001010111: colour_data = 24'b011010101110001101011001;
		13'b0100001011000: colour_data = 24'b001000011000111000100001;
		13'b0100001011001: colour_data = 24'b000110000110110100011000;
		13'b0100001011010: colour_data = 24'b011010101110001101011001;
		13'b0100001011011: colour_data = 24'b011010101110001101011001;
		13'b0100001011100: colour_data = 24'b011010101110001101011001;
		13'b0100001011101: colour_data = 24'b001000011000111000100001;
		13'b0100001011110: colour_data = 24'b001000011000111000100001;
		13'b0100001011111: colour_data = 24'b011010101110001101011001;
		13'b0100001100000: colour_data = 24'b011010101110001101011001;
		13'b0100001100001: colour_data = 24'b001000011000111000100001;
		13'b0100001100010: colour_data = 24'b001000011000111000100001;
		13'b0100001100011: colour_data = 24'b001000011000111000100001;
		13'b0100001100100: colour_data = 24'b011010101110001101011001;
		13'b0100001100101: colour_data = 24'b011010101110001101011001;
		13'b0100001100110: colour_data = 24'b001000011000111000100001;
		13'b0100001100111: colour_data = 24'b000110000110110100011000;
		13'b0100001101000: colour_data = 24'b001000011000111000100001;
		13'b0100001101001: colour_data = 24'b011010101110001101011001;
		13'b0100001101010: colour_data = 24'b011010101110001101011001;
		13'b0100001101011: colour_data = 24'b001000011000111000100001;
		13'b0100001101100: colour_data = 24'b000110000110110100011000;
		13'b0100001101101: colour_data = 24'b011010101110001101011001;
		13'b0100001101110: colour_data = 24'b011010101110001101011001;
		13'b0100001101111: colour_data = 24'b011010101110001101011001;
		13'b0100001110000: colour_data = 24'b001000011000111000100001;
		13'b0100001110001: colour_data = 24'b001000011000111000100001;
		13'b0100001110010: colour_data = 24'b011010101110001101011001;
		13'b0100001110011: colour_data = 24'b011010101110001101011001;
		13'b0100001110100: colour_data = 24'b001000011000111000100001;
		13'b0100001110101: colour_data = 24'b001000011000111000100001;
		13'b0100001110110: colour_data = 24'b001000011000111000100001;
		13'b0100001110111: colour_data = 24'b011010101110001101011001;
		13'b0100001111000: colour_data = 24'b011010101110001101011001;
		13'b0100001111001: colour_data = 24'b001000011000111000100001;
		13'b0100001111010: colour_data = 24'b000110000110110100011000;
		13'b0100001111011: colour_data = 24'b011010101110001101011001;
		13'b0100001111100: colour_data = 24'b011010101110001101011001;
		13'b0100001111101: colour_data = 24'b011010101110001101011001;
		13'b0100001111110: colour_data = 24'b001000011000111000100001;
		13'b0100001111111: colour_data = 24'b000110000110110100011000;
		13'b0100010000000: colour_data = 24'b011010101110001101011001;
		13'b0100010000001: colour_data = 24'b011010101110001101011001;
		13'b0100010000010: colour_data = 24'b011010101110001101011001;
		13'b0100010000011: colour_data = 24'b001000011000111000100001;
		13'b0100010000100: colour_data = 24'b001000011000111000100001;
		13'b0100010000101: colour_data = 24'b011010101110001101011001;
		13'b0100010000110: colour_data = 24'b011010101110001101011001;
		13'b0100010000111: colour_data = 24'b001000011000111000100001;
		13'b0100010001000: colour_data = 24'b000110000110110100011000;
		13'b0100010001001: colour_data = 24'b000110000110110100011000;

		13'b0100100000000: colour_data = 24'b001010101100010100011000;
		13'b0100100000001: colour_data = 24'b011010101110001101011001;
		13'b0100100000010: colour_data = 24'b011010101110001101011001;
		13'b0100100000011: colour_data = 24'b001000011000111000100001;
		13'b0100100000100: colour_data = 24'b001000011000111000100001;
		13'b0100100000101: colour_data = 24'b011010101110001101011001;
		13'b0100100000110: colour_data = 24'b011010101110001101011001;
		13'b0100100000111: colour_data = 24'b001000011000111000100001;
		13'b0100100001000: colour_data = 24'b001000011000111000100001;
		13'b0100100001001: colour_data = 24'b001000011000111000100001;
		13'b0100100001010: colour_data = 24'b011010101110001101011001;
		13'b0100100001011: colour_data = 24'b011010101110001101011001;
		13'b0100100001100: colour_data = 24'b001000011000111000100001;
		13'b0100100001101: colour_data = 24'b000110000110110100011000;
		13'b0100100001110: colour_data = 24'b001000011000111000100001;
		13'b0100100001111: colour_data = 24'b011010101110001101011001;
		13'b0100100010000: colour_data = 24'b011010101110001101011001;
		13'b0100100010001: colour_data = 24'b001000011000111000100001;
		13'b0100100010010: colour_data = 24'b000110000110110100011000;
		13'b0100100010011: colour_data = 24'b011010101110001101011001;
		13'b0100100010100: colour_data = 24'b011010101110001101011001;
		13'b0100100010101: colour_data = 24'b011010101110001101011001;
		13'b0100100010110: colour_data = 24'b001000011000111000100001;
		13'b0100100010111: colour_data = 24'b001000011000111000100001;
		13'b0100100011000: colour_data = 24'b011010101110001101011001;
		13'b0100100011001: colour_data = 24'b011010101110001101011001;
		13'b0100100011010: colour_data = 24'b001000011000111000100001;
		13'b0100100011011: colour_data = 24'b001000011000111000100001;
		13'b0100100011100: colour_data = 24'b001000011000111000100001;
		13'b0100100011101: colour_data = 24'b011010101110001101011001;
		13'b0100100011110: colour_data = 24'b011010101110001101011001;
		13'b0100100011111: colour_data = 24'b001000011000111000100001;
		13'b0100100100000: colour_data = 24'b000110000110110100011000;
		13'b0100100100001: colour_data = 24'b011010101110001101011001;
		13'b0100100100010: colour_data = 24'b011010101110001101011001;
		13'b0100100100011: colour_data = 24'b011010101110001101011001;
		13'b0100100100100: colour_data = 24'b001000011000111000100001;
		13'b0100100100101: colour_data = 24'b000110000110110100011000;
		13'b0100100100110: colour_data = 24'b011010101110001101011001;
		13'b0100100100111: colour_data = 24'b011010101110001101011001;
		13'b0100100101000: colour_data = 24'b011010101110001101011001;
		13'b0100100101001: colour_data = 24'b001000011000111000100001;
		13'b0100100101010: colour_data = 24'b001000011000111000100001;
		13'b0100100101011: colour_data = 24'b011010101110001101011001;
		13'b0100100101100: colour_data = 24'b011010101110001101011001;
		13'b0100100101101: colour_data = 24'b001000011000111000100001;
		13'b0100100101110: colour_data = 24'b001000011000111000100001;
		13'b0100100101111: colour_data = 24'b001000011000111000100001;
		13'b0100100110000: colour_data = 24'b011010101110001101011001;
		13'b0100100110001: colour_data = 24'b011010101110001101011001;
		13'b0100100110010: colour_data = 24'b001000011000111000100001;
		13'b0100100110011: colour_data = 24'b000110000110110100011000;
		13'b0100100110100: colour_data = 24'b001010101100010100011000;
		13'b0100100110101: colour_data = 24'b011010101110001101011001;
		13'b0100100110110: colour_data = 24'b011010101110001101011001;
		13'b0100100110111: colour_data = 24'b001000011000111000100001;
		13'b0100100111000: colour_data = 24'b000110000110110100011000;
		13'b0100100111001: colour_data = 24'b011010101110001101011001;
		13'b0100100111010: colour_data = 24'b011010101110001101011001;
		13'b0100100111011: colour_data = 24'b011010101110001101011001;
		13'b0100100111100: colour_data = 24'b001000011000111000100001;
		13'b0100100111101: colour_data = 24'b001000011000111000100001;
		13'b0100100111110: colour_data = 24'b011010101110001101011001;
		13'b0100100111111: colour_data = 24'b011010101110001101011001;
		13'b0100101000000: colour_data = 24'b001000011000111000100001;
		13'b0100101000001: colour_data = 24'b000110000110110100011000;
		13'b0100101000010: colour_data = 24'b001000011000111000100001;
		13'b0100101000011: colour_data = 24'b011010101110001101011001;
		13'b0100101000100: colour_data = 24'b011010101110001101011001;
		13'b0100101000101: colour_data = 24'b001000011000111000100001;
		13'b0100101000110: colour_data = 24'b000110000110110100011000;
		13'b0100101000111: colour_data = 24'b011010101110001101011001;
		13'b0100101001000: colour_data = 24'b011010101110001101011001;
		13'b0100101001001: colour_data = 24'b011010101110001101011001;
		13'b0100101001010: colour_data = 24'b001000011000111000100001;
		13'b0100101001011: colour_data = 24'b000110000110110100011000;
		13'b0100101001100: colour_data = 24'b011010101110001101011001;
		13'b0100101001101: colour_data = 24'b011010101110001101011001;
		13'b0100101001110: colour_data = 24'b001000011000111000100001;
		13'b0100101001111: colour_data = 24'b001000011000111000100001;
		13'b0100101010000: colour_data = 24'b001000011000111000100001;
		13'b0100101010001: colour_data = 24'b011010101110001101011001;
		13'b0100101010010: colour_data = 24'b011010101110001101011001;
		13'b0100101010011: colour_data = 24'b001000011000111000100001;
		13'b0100101010100: colour_data = 24'b000110000110110100011000;
		13'b0100101010101: colour_data = 24'b001000011000111000100001;
		13'b0100101010110: colour_data = 24'b011010101110001101011001;
		13'b0100101010111: colour_data = 24'b011010101110001101011001;
		13'b0100101011000: colour_data = 24'b001000011000111000100001;
		13'b0100101011001: colour_data = 24'b000110000110110100011000;
		13'b0100101011010: colour_data = 24'b011010101110001101011001;
		13'b0100101011011: colour_data = 24'b011010101110001101011001;
		13'b0100101011100: colour_data = 24'b011010101110001101011001;
		13'b0100101011101: colour_data = 24'b001000011000111000100001;
		13'b0100101011110: colour_data = 24'b001000011000111000100001;
		13'b0100101011111: colour_data = 24'b011010101110001101011001;
		13'b0100101100000: colour_data = 24'b011010101110001101011001;
		13'b0100101100001: colour_data = 24'b001000011000111000100001;
		13'b0100101100010: colour_data = 24'b001000011000111000100001;
		13'b0100101100011: colour_data = 24'b001000011000111000100001;
		13'b0100101100100: colour_data = 24'b011010101110001101011001;
		13'b0100101100101: colour_data = 24'b011010101110001101011001;
		13'b0100101100110: colour_data = 24'b001000011000111000100001;
		13'b0100101100111: colour_data = 24'b000110000110110100011000;
		13'b0100101101000: colour_data = 24'b001000011000111000100001;
		13'b0100101101001: colour_data = 24'b011010101110001101011001;
		13'b0100101101010: colour_data = 24'b011010101110001101011001;
		13'b0100101101011: colour_data = 24'b001000011000111000100001;
		13'b0100101101100: colour_data = 24'b000110000110110100011000;
		13'b0100101101101: colour_data = 24'b011010101110001101011001;
		13'b0100101101110: colour_data = 24'b011010101110001101011001;
		13'b0100101101111: colour_data = 24'b011010101110001101011001;
		13'b0100101110000: colour_data = 24'b001000011000111000100001;
		13'b0100101110001: colour_data = 24'b001000011000111000100001;
		13'b0100101110010: colour_data = 24'b011010101110001101011001;
		13'b0100101110011: colour_data = 24'b011010101110001101011001;
		13'b0100101110100: colour_data = 24'b001000011000111000100001;
		13'b0100101110101: colour_data = 24'b001000011000111000100001;
		13'b0100101110110: colour_data = 24'b001000011000111000100001;
		13'b0100101110111: colour_data = 24'b011010101110001101011001;
		13'b0100101111000: colour_data = 24'b011010101110001101011001;
		13'b0100101111001: colour_data = 24'b001000011000111000100001;
		13'b0100101111010: colour_data = 24'b000110000110110100011000;
		13'b0100101111011: colour_data = 24'b011010101110001101011001;
		13'b0100101111100: colour_data = 24'b011010101110001101011001;
		13'b0100101111101: colour_data = 24'b011010101110001101011001;
		13'b0100101111110: colour_data = 24'b001000011000111000100001;
		13'b0100101111111: colour_data = 24'b000110000110110100011000;
		13'b0100110000000: colour_data = 24'b011010101110001101011001;
		13'b0100110000001: colour_data = 24'b011010101110001101011001;
		13'b0100110000010: colour_data = 24'b011010101110001101011001;
		13'b0100110000011: colour_data = 24'b001000011000111000100001;
		13'b0100110000100: colour_data = 24'b001000011000111000100001;
		13'b0100110000101: colour_data = 24'b011010101110001101011001;
		13'b0100110000110: colour_data = 24'b011010101110001101011001;
		13'b0100110000111: colour_data = 24'b001000011000111000100001;
		13'b0100110001000: colour_data = 24'b000110000110110100011000;
		13'b0100110001001: colour_data = 24'b000110000110110100011000;

		13'b0101000000000: colour_data = 24'b001010101100010100011000;
		13'b0101000000001: colour_data = 24'b011010101110001101011001;
		13'b0101000000010: colour_data = 24'b011010101110001101011001;
		13'b0101000000011: colour_data = 24'b001000011000111000100001;
		13'b0101000000100: colour_data = 24'b001000011000111000100001;
		13'b0101000000101: colour_data = 24'b011010101110001101011001;
		13'b0101000000110: colour_data = 24'b011010101110001101011001;
		13'b0101000000111: colour_data = 24'b000110000110110100011000;
		13'b0101000001000: colour_data = 24'b001000011000111000100001;
		13'b0101000001001: colour_data = 24'b000110000110110100011000;
		13'b0101000001010: colour_data = 24'b011010101110001101011001;
		13'b0101000001011: colour_data = 24'b011010101110001101011001;
		13'b0101000001100: colour_data = 24'b000110000110110100011000;
		13'b0101000001101: colour_data = 24'b000110000110110100011000;
		13'b0101000001110: colour_data = 24'b001000011000111000100001;
		13'b0101000001111: colour_data = 24'b011010101110001101011001;
		13'b0101000010000: colour_data = 24'b011010101110001101011001;
		13'b0101000010001: colour_data = 24'b001000011000111000100001;
		13'b0101000010010: colour_data = 24'b000110000110110100011000;
		13'b0101000010011: colour_data = 24'b011010101110001101011001;
		13'b0101000010100: colour_data = 24'b011010101110001101011001;
		13'b0101000010101: colour_data = 24'b011010101110001101011001;
		13'b0101000010110: colour_data = 24'b001000011000111000100001;
		13'b0101000010111: colour_data = 24'b000110000110110100011000;
		13'b0101000011000: colour_data = 24'b001010101100010100011000;
		13'b0101000011001: colour_data = 24'b011010101110001101011001;
		13'b0101000011010: colour_data = 24'b000110000110110100011000;
		13'b0101000011011: colour_data = 24'b001000011000111000100001;
		13'b0101000011100: colour_data = 24'b001000011000111000100001;
		13'b0101000011101: colour_data = 24'b011010101110001101011001;
		13'b0101000011110: colour_data = 24'b011010101110001101011001;
		13'b0101000011111: colour_data = 24'b000110000110110100011000;
		13'b0101000100000: colour_data = 24'b000110000110110100011000;
		13'b0101000100001: colour_data = 24'b001010101100010100011000;
		13'b0101000100010: colour_data = 24'b011010101110001101011001;
		13'b0101000100011: colour_data = 24'b011010101110001101011001;
		13'b0101000100100: colour_data = 24'b001000011000111000100001;
		13'b0101000100101: colour_data = 24'b000110000110110100011000;
		13'b0101000100110: colour_data = 24'b011010101110001101011001;
		13'b0101000100111: colour_data = 24'b011010101110001101011001;
		13'b0101000101000: colour_data = 24'b011010101110001101011001;
		13'b0101000101001: colour_data = 24'b001000011000111000100001;
		13'b0101000101010: colour_data = 24'b000110000110110100011000;
		13'b0101000101011: colour_data = 24'b001010101100010100011000;
		13'b0101000101100: colour_data = 24'b011010101110001101011001;
		13'b0101000101101: colour_data = 24'b000110000110110100011000;
		13'b0101000101110: colour_data = 24'b001000011000111000100001;
		13'b0101000101111: colour_data = 24'b001000011000111000100001;
		13'b0101000110000: colour_data = 24'b011010101110001101011001;
		13'b0101000110001: colour_data = 24'b011010101110001101011001;
		13'b0101000110010: colour_data = 24'b000110000110110100011000;
		13'b0101000110011: colour_data = 24'b000110000110110100011000;
		13'b0101000110100: colour_data = 24'b001010101100010100011000;
		13'b0101000110101: colour_data = 24'b011010101110001101011001;
		13'b0101000110110: colour_data = 24'b011010101110001101011001;
		13'b0101000110111: colour_data = 24'b001000011000111000100001;
		13'b0101000111000: colour_data = 24'b000110000110110100011000;
		13'b0101000111001: colour_data = 24'b011010101110001101011001;
		13'b0101000111010: colour_data = 24'b011010101110001101011001;
		13'b0101000111011: colour_data = 24'b011010101110001101011001;
		13'b0101000111100: colour_data = 24'b001000011000111000100001;
		13'b0101000111101: colour_data = 24'b000110000110110100011000;
		13'b0101000111110: colour_data = 24'b011010101110001101011001;
		13'b0101000111111: colour_data = 24'b011010101110001101011001;
		13'b0101001000000: colour_data = 24'b000110000110110100011000;
		13'b0101001000001: colour_data = 24'b000110000110110100011000;
		13'b0101001000010: colour_data = 24'b001000011000111000100001;
		13'b0101001000011: colour_data = 24'b011010101110001101011001;
		13'b0101001000100: colour_data = 24'b011010101110001101011001;
		13'b0101001000101: colour_data = 24'b000110000110110100011000;
		13'b0101001000110: colour_data = 24'b000110000110110100011000;
		13'b0101001000111: colour_data = 24'b011010101110001101011001;
		13'b0101001001000: colour_data = 24'b011010101110001101011001;
		13'b0101001001001: colour_data = 24'b011010101110001101011001;
		13'b0101001001010: colour_data = 24'b001000011000111000100001;
		13'b0101001001011: colour_data = 24'b000110000110110100011000;
		13'b0101001001100: colour_data = 24'b001010101100010100011000;
		13'b0101001001101: colour_data = 24'b011010101110001101011001;
		13'b0101001001110: colour_data = 24'b000110000110110100011000;
		13'b0101001001111: colour_data = 24'b001000011000111000100001;
		13'b0101001010000: colour_data = 24'b001000011000111000100001;
		13'b0101001010001: colour_data = 24'b011010101110001101011001;
		13'b0101001010010: colour_data = 24'b011010101110001101011001;
		13'b0101001010011: colour_data = 24'b000110000110110100011000;
		13'b0101001010100: colour_data = 24'b000110000110110100011000;
		13'b0101001010101: colour_data = 24'b000110000110110100011000;
		13'b0101001010110: colour_data = 24'b011010101110001101011001;
		13'b0101001010111: colour_data = 24'b011010101110001101011001;
		13'b0101001011000: colour_data = 24'b000110000110110100011000;
		13'b0101001011001: colour_data = 24'b000110000110110100011000;
		13'b0101001011010: colour_data = 24'b011010101110001101011001;
		13'b0101001011011: colour_data = 24'b011010101110001101011001;
		13'b0101001011100: colour_data = 24'b011010101110001101011001;
		13'b0101001011101: colour_data = 24'b001000011000111000100001;
		13'b0101001011110: colour_data = 24'b000110000110110100011000;
		13'b0101001011111: colour_data = 24'b001010101100010100011000;
		13'b0101001100000: colour_data = 24'b011010101110001101011001;
		13'b0101001100001: colour_data = 24'b000110000110110100011000;
		13'b0101001100010: colour_data = 24'b001000011000111000100001;
		13'b0101001100011: colour_data = 24'b001000011000111000100001;
		13'b0101001100100: colour_data = 24'b011010101110001101011001;
		13'b0101001100101: colour_data = 24'b011010101110001101011001;
		13'b0101001100110: colour_data = 24'b000110000110110100011000;
		13'b0101001100111: colour_data = 24'b000110000110110100011000;
		13'b0101001101000: colour_data = 24'b000110000110110100011000;
		13'b0101001101001: colour_data = 24'b011010101110001101011001;
		13'b0101001101010: colour_data = 24'b011010101110001101011001;
		13'b0101001101011: colour_data = 24'b001000011000111000100001;
		13'b0101001101100: colour_data = 24'b000110000110110100011000;
		13'b0101001101101: colour_data = 24'b011010101110001101011001;
		13'b0101001101110: colour_data = 24'b011010101110001101011001;
		13'b0101001101111: colour_data = 24'b011010101110001101011001;
		13'b0101001110000: colour_data = 24'b001000011000111000100001;
		13'b0101001110001: colour_data = 24'b000110000110110100011000;
		13'b0101001110010: colour_data = 24'b001010101100010100011000;
		13'b0101001110011: colour_data = 24'b011010101110001101011001;
		13'b0101001110100: colour_data = 24'b000110000110110100011000;
		13'b0101001110101: colour_data = 24'b001000011000111000100001;
		13'b0101001110110: colour_data = 24'b001000011000111000100001;
		13'b0101001110111: colour_data = 24'b011010101110001101011001;
		13'b0101001111000: colour_data = 24'b011010101110001101011001;
		13'b0101001111001: colour_data = 24'b000110000110110100011000;
		13'b0101001111010: colour_data = 24'b000110000110110100011000;
		13'b0101001111011: colour_data = 24'b011010101110001101011001;
		13'b0101001111100: colour_data = 24'b011010101110001101011001;
		13'b0101001111101: colour_data = 24'b011010101110001101011001;
		13'b0101001111110: colour_data = 24'b001000011000111000100001;
		13'b0101001111111: colour_data = 24'b000110000110110100011000;
		13'b0101010000000: colour_data = 24'b001010101100010100011000;
		13'b0101010000001: colour_data = 24'b011010101110001101011001;
		13'b0101010000010: colour_data = 24'b011010101110001101011001;
		13'b0101010000011: colour_data = 24'b001000011000111000100001;
		13'b0101010000100: colour_data = 24'b001000011000111000100001;
		13'b0101010000101: colour_data = 24'b011010101110001101011001;
		13'b0101010000110: colour_data = 24'b011010101110001101011001;
		13'b0101010000111: colour_data = 24'b000110000110110100011000;
		13'b0101010001000: colour_data = 24'b000110000110110100011000;
		13'b0101010001001: colour_data = 24'b000110000110110100011000;

		13'b0101100000000: colour_data = 24'b111111110000000010010110;
		13'b0101100000001: colour_data = 24'b001010101100010100011000;
		13'b0101100000010: colour_data = 24'b011010101110001101011001;
		13'b0101100000011: colour_data = 24'b000110000110110100011000;
		13'b0101100000100: colour_data = 24'b000110000110110100011000;
		13'b0101100000101: colour_data = 24'b011010101110001101011001;
		13'b0101100000110: colour_data = 24'b011010101110001101011001;
		13'b0101100000111: colour_data = 24'b000110000110110100011000;
		13'b0101100001000: colour_data = 24'b000110000110110100011000;
		13'b0101100001001: colour_data = 24'b001000011000111000100001;
		13'b0101100001010: colour_data = 24'b001010101100010100011000;
		13'b0101100001011: colour_data = 24'b011010101110001101011001;
		13'b0101100001100: colour_data = 24'b000110000110110100011000;
		13'b0101100001101: colour_data = 24'b000110000110110100011000;
		13'b0101100001110: colour_data = 24'b000110000110110100011000;
		13'b0101100001111: colour_data = 24'b011010101110001101011001;
		13'b0101100010000: colour_data = 24'b011010101110001101011001;
		13'b0101100010001: colour_data = 24'b000110000110110100011000;
		13'b0101100010010: colour_data = 24'b000110000110110100011000;
		13'b0101100010011: colour_data = 24'b011010101110001101011001;
		13'b0101100010100: colour_data = 24'b011010101110001101011001;
		13'b0101100010101: colour_data = 24'b011010101110001101011001;
		13'b0101100010110: colour_data = 24'b000110000110110100011000;
		13'b0101100010111: colour_data = 24'b001000011000111000100001;
		13'b0101100011000: colour_data = 24'b000110000110110100011000;
		13'b0101100011001: colour_data = 24'b011010101110001101011001;
		13'b0101100011010: colour_data = 24'b000110000110110100011000;
		13'b0101100011011: colour_data = 24'b000110000110110100011000;
		13'b0101100011100: colour_data = 24'b000110000110110100011000;
		13'b0101100011101: colour_data = 24'b011010101110001101011001;
		13'b0101100011110: colour_data = 24'b011010101110001101011001;
		13'b0101100011111: colour_data = 24'b000110000110110100011000;
		13'b0101100100000: colour_data = 24'b000110000110110100011000;
		13'b0101100100001: colour_data = 24'b000110000110110100011000;
		13'b0101100100010: colour_data = 24'b001010101100010100011000;
		13'b0101100100011: colour_data = 24'b011010101110001101011001;
		13'b0101100100100: colour_data = 24'b000110000110110100011000;
		13'b0101100100101: colour_data = 24'b000110000110110100011000;
		13'b0101100100110: colour_data = 24'b011010101110001101011001;
		13'b0101100100111: colour_data = 24'b011010101110001101011001;
		13'b0101100101000: colour_data = 24'b011010101110001101011001;
		13'b0101100101001: colour_data = 24'b000110000110110100011000;
		13'b0101100101010: colour_data = 24'b001000011000111000100001;
		13'b0101100101011: colour_data = 24'b000110000110110100011000;
		13'b0101100101100: colour_data = 24'b011010101110001101011001;
		13'b0101100101101: colour_data = 24'b000110000110110100011000;
		13'b0101100101110: colour_data = 24'b000110000110110100011000;
		13'b0101100101111: colour_data = 24'b000110000110110100011000;
		13'b0101100110000: colour_data = 24'b011010101110001101011001;
		13'b0101100110001: colour_data = 24'b011010101110001101011001;
		13'b0101100110010: colour_data = 24'b000110000110110100011000;
		13'b0101100110011: colour_data = 24'b000110000110110100011000;
		13'b0101100110100: colour_data = 24'b000110000110110100011000;
		13'b0101100110101: colour_data = 24'b001010101100010100011000;
		13'b0101100110110: colour_data = 24'b011010101110001101011001;
		13'b0101100110111: colour_data = 24'b000110000110110100011000;
		13'b0101100111000: colour_data = 24'b000110000110110100011000;
		13'b0101100111001: colour_data = 24'b011010101110001101011001;
		13'b0101100111010: colour_data = 24'b011010101110001101011001;
		13'b0101100111011: colour_data = 24'b011010101110001101011001;
		13'b0101100111100: colour_data = 24'b000110000110110100011000;
		13'b0101100111101: colour_data = 24'b001000011000111000100001;
		13'b0101100111110: colour_data = 24'b001010101100010100011000;
		13'b0101100111111: colour_data = 24'b011010101110001101011001;
		13'b0101101000000: colour_data = 24'b000110000110110100011000;
		13'b0101101000001: colour_data = 24'b000110000110110100011000;
		13'b0101101000010: colour_data = 24'b000110000110110100011000;
		13'b0101101000011: colour_data = 24'b011010101110001101011001;
		13'b0101101000100: colour_data = 24'b011010101110001101011001;
		13'b0101101000101: colour_data = 24'b000110000110110100011000;
		13'b0101101000110: colour_data = 24'b000110000110110100011000;
		13'b0101101000111: colour_data = 24'b011010101110001101011001;
		13'b0101101001000: colour_data = 24'b011010101110001101011001;
		13'b0101101001001: colour_data = 24'b011010101110001101011001;
		13'b0101101001010: colour_data = 24'b000110000110110100011000;
		13'b0101101001011: colour_data = 24'b000110000110110100011000;
		13'b0101101001100: colour_data = 24'b000110000110110100011000;
		13'b0101101001101: colour_data = 24'b011010101110001101011001;
		13'b0101101001110: colour_data = 24'b000110000110110100011000;
		13'b0101101001111: colour_data = 24'b000110000110110100011000;
		13'b0101101010000: colour_data = 24'b000110000110110100011000;
		13'b0101101010001: colour_data = 24'b011010101110001101011001;
		13'b0101101010010: colour_data = 24'b011010101110001101011001;
		13'b0101101010011: colour_data = 24'b000110000110110100011000;
		13'b0101101010100: colour_data = 24'b000110000110110100011000;
		13'b0101101010101: colour_data = 24'b001000011000111000100001;
		13'b0101101010110: colour_data = 24'b001010101100010100011000;
		13'b0101101010111: colour_data = 24'b011010101110001101011001;
		13'b0101101011000: colour_data = 24'b000110000110110100011000;
		13'b0101101011001: colour_data = 24'b000110000110110100011000;
		13'b0101101011010: colour_data = 24'b011010101110001101011001;
		13'b0101101011011: colour_data = 24'b011010101110001101011001;
		13'b0101101011100: colour_data = 24'b011010101110001101011001;
		13'b0101101011101: colour_data = 24'b000110000110110100011000;
		13'b0101101011110: colour_data = 24'b001000011000111000100001;
		13'b0101101011111: colour_data = 24'b000110000110110100011000;
		13'b0101101100000: colour_data = 24'b011010101110001101011001;
		13'b0101101100001: colour_data = 24'b000110000110110100011000;
		13'b0101101100010: colour_data = 24'b000110000110110100011000;
		13'b0101101100011: colour_data = 24'b000110000110110100011000;
		13'b0101101100100: colour_data = 24'b011010101110001101011001;
		13'b0101101100101: colour_data = 24'b011010101110001101011001;
		13'b0101101100110: colour_data = 24'b000110000110110100011000;
		13'b0101101100111: colour_data = 24'b000110000110110100011000;
		13'b0101101101000: colour_data = 24'b001000011000111000100001;
		13'b0101101101001: colour_data = 24'b001010101100010100011000;
		13'b0101101101010: colour_data = 24'b011010101110001101011001;
		13'b0101101101011: colour_data = 24'b000110000110110100011000;
		13'b0101101101100: colour_data = 24'b000110000110110100011000;
		13'b0101101101101: colour_data = 24'b011010101110001101011001;
		13'b0101101101110: colour_data = 24'b011010101110001101011001;
		13'b0101101101111: colour_data = 24'b011010101110001101011001;
		13'b0101101110000: colour_data = 24'b000110000110110100011000;
		13'b0101101110001: colour_data = 24'b001000011000111000100001;
		13'b0101101110010: colour_data = 24'b000110000110110100011000;
		13'b0101101110011: colour_data = 24'b011010101110001101011001;
		13'b0101101110100: colour_data = 24'b000110000110110100011000;
		13'b0101101110101: colour_data = 24'b000110000110110100011000;
		13'b0101101110110: colour_data = 24'b000110000110110100011000;
		13'b0101101110111: colour_data = 24'b001010101100010100011000;
		13'b0101101111000: colour_data = 24'b011010101110001101011001;
		13'b0101101111001: colour_data = 24'b000110000110110100011000;
		13'b0101101111010: colour_data = 24'b000110000110110100011000;
		13'b0101101111011: colour_data = 24'b011010101110001101011001;
		13'b0101101111100: colour_data = 24'b011010101110001101011001;
		13'b0101101111101: colour_data = 24'b011010101110001101011001;
		13'b0101101111110: colour_data = 24'b000110000110110100011000;
		13'b0101101111111: colour_data = 24'b000110000110110100011000;
		13'b0101110000000: colour_data = 24'b000110000110110100011000;
		13'b0101110000001: colour_data = 24'b011010101110001101011001;
		13'b0101110000010: colour_data = 24'b011010101110001101011001;
		13'b0101110000011: colour_data = 24'b000110000110110100011000;
		13'b0101110000100: colour_data = 24'b000110000110110100011000;
		13'b0101110000101: colour_data = 24'b011010101110001101011001;
		13'b0101110000110: colour_data = 24'b011010101110001101011001;
		13'b0101110000111: colour_data = 24'b000110000110110100011000;
		13'b0101110001000: colour_data = 24'b000110000110110100011000;
		13'b0101110001001: colour_data = 24'b111111110000000010010110;

		13'b0110000000000: colour_data = 24'b111111110000000010010110;
		13'b0110000000001: colour_data = 24'b111111110000000010010110;
		13'b0110000000010: colour_data = 24'b011010101110001101011001;
		13'b0110000000011: colour_data = 24'b000110000110110100011000;
		13'b0110000000100: colour_data = 24'b000110000110110100011000;
		13'b0110000000101: colour_data = 24'b011010101110001101011001;
		13'b0110000000110: colour_data = 24'b011010101110001101011001;
		13'b0110000000111: colour_data = 24'b000110000110110100011000;
		13'b0110000001000: colour_data = 24'b000110000110110100011000;
		13'b0110000001001: colour_data = 24'b001000011000111000100001;
		13'b0110000001010: colour_data = 24'b000110000101000100011000;
		13'b0110000001011: colour_data = 24'b001010101100010100011000;
		13'b0110000001100: colour_data = 24'b000110000110110100011000;
		13'b0110000001101: colour_data = 24'b000110000110110100011000;
		13'b0110000001110: colour_data = 24'b000110000110110100011000;
		13'b0110000001111: colour_data = 24'b011010101110001101011001;
		13'b0110000010000: colour_data = 24'b011010101110001101011001;
		13'b0110000010001: colour_data = 24'b000110000110110100011000;
		13'b0110000010010: colour_data = 24'b001000011000111000100001;
		13'b0110000010011: colour_data = 24'b011010101110001101011001;
		13'b0110000010100: colour_data = 24'b011010101110001101011001;
		13'b0110000010101: colour_data = 24'b011010101110001101011001;
		13'b0110000010110: colour_data = 24'b000110000110110100011000;
		13'b0110000010111: colour_data = 24'b001000011000111000100001;
		13'b0110000011000: colour_data = 24'b000110000110110100011000;
		13'b0110000011001: colour_data = 24'b001010101100010100011000;
		13'b0110000011010: colour_data = 24'b000110000110110100011000;
		13'b0110000011011: colour_data = 24'b000110000110110100011000;
		13'b0110000011100: colour_data = 24'b000110000110110100011000;
		13'b0110000011101: colour_data = 24'b011010101110001101011001;
		13'b0110000011110: colour_data = 24'b011010101110001101011001;
		13'b0110000011111: colour_data = 24'b000110000110110100011000;
		13'b0110000100000: colour_data = 24'b001000011000111000100001;
		13'b0110000100001: colour_data = 24'b000110000110110100011000;
		13'b0110000100010: colour_data = 24'b000110000101000100011000;
		13'b0110000100011: colour_data = 24'b011010101110001101011001;
		13'b0110000100100: colour_data = 24'b000110000110110100011000;
		13'b0110000100101: colour_data = 24'b000110000110110100011000;
		13'b0110000100110: colour_data = 24'b011010101110001101011001;
		13'b0110000100111: colour_data = 24'b011010101110001101011001;
		13'b0110000101000: colour_data = 24'b011010101110001101011001;
		13'b0110000101001: colour_data = 24'b000110000110110100011000;
		13'b0110000101010: colour_data = 24'b001000011000111000100001;
		13'b0110000101011: colour_data = 24'b000110000110110100011000;
		13'b0110000101100: colour_data = 24'b001010101100010100011000;
		13'b0110000101101: colour_data = 24'b000110000110110100011000;
		13'b0110000101110: colour_data = 24'b000110000110110100011000;
		13'b0110000101111: colour_data = 24'b000110000110110100011000;
		13'b0110000110000: colour_data = 24'b011010101110001101011001;
		13'b0110000110001: colour_data = 24'b011010101110001101011001;
		13'b0110000110010: colour_data = 24'b000110000110110100011000;
		13'b0110000110011: colour_data = 24'b001000011000111000100001;
		13'b0110000110100: colour_data = 24'b000110000110110100011000;
		13'b0110000110101: colour_data = 24'b000110000101000100011000;
		13'b0110000110110: colour_data = 24'b011010101110001101011001;
		13'b0110000110111: colour_data = 24'b000110000110110100011000;
		13'b0110000111000: colour_data = 24'b000110000110110100011000;
		13'b0110000111001: colour_data = 24'b011010101110001101011001;
		13'b0110000111010: colour_data = 24'b011010101110001101011001;
		13'b0110000111011: colour_data = 24'b011010101110001101011001;
		13'b0110000111100: colour_data = 24'b000110000110110100011000;
		13'b0110000111101: colour_data = 24'b001000011000111000100001;
		13'b0110000111110: colour_data = 24'b000110000101000100011000;
		13'b0110000111111: colour_data = 24'b001010101100010100011000;
		13'b0110001000000: colour_data = 24'b000110000110110100011000;
		13'b0110001000001: colour_data = 24'b000110000110110100011000;
		13'b0110001000010: colour_data = 24'b000110000110110100011000;
		13'b0110001000011: colour_data = 24'b011010101110001101011001;
		13'b0110001000100: colour_data = 24'b011010101110001101011001;
		13'b0110001000101: colour_data = 24'b000110000110110100011000;
		13'b0110001000110: colour_data = 24'b001000011000111000100001;
		13'b0110001000111: colour_data = 24'b011010101110001101011001;
		13'b0110001001000: colour_data = 24'b011010101110001101011001;
		13'b0110001001001: colour_data = 24'b011010101110001101011001;
		13'b0110001001010: colour_data = 24'b000110000110110100011000;
		13'b0110001001011: colour_data = 24'b001000011000111000100001;
		13'b0110001001100: colour_data = 24'b000110000110110100011000;
		13'b0110001001101: colour_data = 24'b001010101100010100011000;
		13'b0110001001110: colour_data = 24'b000110000110110100011000;
		13'b0110001001111: colour_data = 24'b000110000110110100011000;
		13'b0110001010000: colour_data = 24'b000110000110110100011000;
		13'b0110001010001: colour_data = 24'b011010101110001101011001;
		13'b0110001010010: colour_data = 24'b011010101110001101011001;
		13'b0110001010011: colour_data = 24'b000110000110110100011000;
		13'b0110001010100: colour_data = 24'b001000011000111000100001;
		13'b0110001010101: colour_data = 24'b001000011000111000100001;
		13'b0110001010110: colour_data = 24'b000110000101000100011000;
		13'b0110001010111: colour_data = 24'b011010101110001101011001;
		13'b0110001011000: colour_data = 24'b000110000110110100011000;
		13'b0110001011001: colour_data = 24'b000110000110110100011000;
		13'b0110001011010: colour_data = 24'b011010101110001101011001;
		13'b0110001011011: colour_data = 24'b011010101110001101011001;
		13'b0110001011100: colour_data = 24'b011010101110001101011001;
		13'b0110001011101: colour_data = 24'b000110000110110100011000;
		13'b0110001011110: colour_data = 24'b001000011000111000100001;
		13'b0110001011111: colour_data = 24'b000110000110110100011000;
		13'b0110001100000: colour_data = 24'b001010101100010100011000;
		13'b0110001100001: colour_data = 24'b000110000110110100011000;
		13'b0110001100010: colour_data = 24'b000110000110110100011000;
		13'b0110001100011: colour_data = 24'b000110000110110100011000;
		13'b0110001100100: colour_data = 24'b011010101110001101011001;
		13'b0110001100101: colour_data = 24'b011010101110001101011001;
		13'b0110001100110: colour_data = 24'b000110000110110100011000;
		13'b0110001100111: colour_data = 24'b001000011000111000100001;
		13'b0110001101000: colour_data = 24'b001000011000111000100001;
		13'b0110001101001: colour_data = 24'b000110000101000100011000;
		13'b0110001101010: colour_data = 24'b011010101110001101011001;
		13'b0110001101011: colour_data = 24'b000110000110110100011000;
		13'b0110001101100: colour_data = 24'b000110000110110100011000;
		13'b0110001101101: colour_data = 24'b011010101110001101011001;
		13'b0110001101110: colour_data = 24'b011010101110001101011001;
		13'b0110001101111: colour_data = 24'b011010101110001101011001;
		13'b0110001110000: colour_data = 24'b000110000110110100011000;
		13'b0110001110001: colour_data = 24'b001000011000111000100001;
		13'b0110001110010: colour_data = 24'b000110000110110100011000;
		13'b0110001110011: colour_data = 24'b001010101100010100011000;
		13'b0110001110100: colour_data = 24'b000110000110110100011000;
		13'b0110001110101: colour_data = 24'b000110000110110100011000;
		13'b0110001110110: colour_data = 24'b000110000110110100011000;
		13'b0110001110111: colour_data = 24'b000110000101000100011000;
		13'b0110001111000: colour_data = 24'b001010101100010100011000;
		13'b0110001111001: colour_data = 24'b000110000110110100011000;
		13'b0110001111010: colour_data = 24'b000110000110110100011000;
		13'b0110001111011: colour_data = 24'b011010101110001101011001;
		13'b0110001111100: colour_data = 24'b011010101110001101011001;
		13'b0110001111101: colour_data = 24'b011010101110001101011001;
		13'b0110001111110: colour_data = 24'b000110000110110100011000;
		13'b0110001111111: colour_data = 24'b001000011000111000100001;
		13'b0110010000000: colour_data = 24'b000110000110110100011000;
		13'b0110010000001: colour_data = 24'b001010101100010100011000;
		13'b0110010000010: colour_data = 24'b011010101110001101011001;
		13'b0110010000011: colour_data = 24'b000110000110110100011000;
		13'b0110010000100: colour_data = 24'b000110000110110100011000;
		13'b0110010000101: colour_data = 24'b011010101110001101011001;
		13'b0110010000110: colour_data = 24'b011010101110001101011001;
		13'b0110010000111: colour_data = 24'b000110000110110100011000;
		13'b0110010001000: colour_data = 24'b111111110000000010010110;
		13'b0110010001001: colour_data = 24'b111111110000000010010110;

		13'b0110100000000: colour_data = 24'b111111110000000010010110;
		13'b0110100000001: colour_data = 24'b111111110000000010010110;
		13'b0110100000010: colour_data = 24'b001010101100010100011000;
		13'b0110100000011: colour_data = 24'b000110000110110100011000;
		13'b0110100000100: colour_data = 24'b000110000110110100011000;
		13'b0110100000101: colour_data = 24'b011010101110001101011001;
		13'b0110100000110: colour_data = 24'b011010101110001101011001;
		13'b0110100000111: colour_data = 24'b000110000110110100011000;
		13'b0110100001000: colour_data = 24'b001000011000111000100001;
		13'b0110100001001: colour_data = 24'b001000011000111000100001;
		13'b0110100001010: colour_data = 24'b000110000101000100011000;
		13'b0110100001011: colour_data = 24'b000110000110110100011000;
		13'b0110100001100: colour_data = 24'b000110000110110100011000;
		13'b0110100001101: colour_data = 24'b000110000110110100011000;
		13'b0110100001110: colour_data = 24'b000110000110110100011000;
		13'b0110100001111: colour_data = 24'b011010101110001101011001;
		13'b0110100010000: colour_data = 24'b011010101110001101011001;
		13'b0110100010001: colour_data = 24'b001000011000111000100001;
		13'b0110100010010: colour_data = 24'b001000011000111000100001;
		13'b0110100010011: colour_data = 24'b011010101110001101011001;
		13'b0110100010100: colour_data = 24'b011010101110001101011001;
		13'b0110100010101: colour_data = 24'b011010101110001101011001;
		13'b0110100010110: colour_data = 24'b001000011000111000100001;
		13'b0110100010111: colour_data = 24'b001000011000111000100001;
		13'b0110100011000: colour_data = 24'b000110000110110100011000;
		13'b0110100011001: colour_data = 24'b000110000110110100011000;
		13'b0110100011010: colour_data = 24'b000110000110110100011000;
		13'b0110100011011: colour_data = 24'b000110000110110100011000;
		13'b0110100011100: colour_data = 24'b000110000110110100011000;
		13'b0110100011101: colour_data = 24'b011010101110001101011001;
		13'b0110100011110: colour_data = 24'b011010101110001101011001;
		13'b0110100011111: colour_data = 24'b000110000110110100011000;
		13'b0110100100000: colour_data = 24'b001000011000111000100001;
		13'b0110100100001: colour_data = 24'b000110000110110100011000;
		13'b0110100100010: colour_data = 24'b000110000101000100011000;
		13'b0110100100011: colour_data = 24'b001010101100010100011000;
		13'b0110100100100: colour_data = 24'b000110000110110100011000;
		13'b0110100100101: colour_data = 24'b000110000110110100011000;
		13'b0110100100110: colour_data = 24'b011010101110001101011001;
		13'b0110100100111: colour_data = 24'b011010101110001101011001;
		13'b0110100101000: colour_data = 24'b011010101110001101011001;
		13'b0110100101001: colour_data = 24'b001000011000111000100001;
		13'b0110100101010: colour_data = 24'b001000011000111000100001;
		13'b0110100101011: colour_data = 24'b000110000110110100011000;
		13'b0110100101100: colour_data = 24'b000110000110110100011000;
		13'b0110100101101: colour_data = 24'b000110000110110100011000;
		13'b0110100101110: colour_data = 24'b000110000110110100011000;
		13'b0110100101111: colour_data = 24'b000110000110110100011000;
		13'b0110100110000: colour_data = 24'b011010101110001101011001;
		13'b0110100110001: colour_data = 24'b011010101110001101011001;
		13'b0110100110010: colour_data = 24'b000110000110110100011000;
		13'b0110100110011: colour_data = 24'b001000011000111000100001;
		13'b0110100110100: colour_data = 24'b000110000110110100011000;
		13'b0110100110101: colour_data = 24'b000110000101000100011000;
		13'b0110100110110: colour_data = 24'b001010101100010100011000;
		13'b0110100110111: colour_data = 24'b000110000110110100011000;
		13'b0110100111000: colour_data = 24'b000110000110110100011000;
		13'b0110100111001: colour_data = 24'b011010101110001101011001;
		13'b0110100111010: colour_data = 24'b011010101110001101011001;
		13'b0110100111011: colour_data = 24'b011010101110001101011001;
		13'b0110100111100: colour_data = 24'b001000011000111000100001;
		13'b0110100111101: colour_data = 24'b001000011000111000100001;
		13'b0110100111110: colour_data = 24'b000110000101000100011000;
		13'b0110100111111: colour_data = 24'b000110000110110100011000;
		13'b0110101000000: colour_data = 24'b000110000110110100011000;
		13'b0110101000001: colour_data = 24'b000110000110110100011000;
		13'b0110101000010: colour_data = 24'b000110000110110100011000;
		13'b0110101000011: colour_data = 24'b011010101110001101011001;
		13'b0110101000100: colour_data = 24'b011010101110001101011001;
		13'b0110101000101: colour_data = 24'b000110000110110100011000;
		13'b0110101000110: colour_data = 24'b001000011000111000100001;
		13'b0110101000111: colour_data = 24'b011010101110001101011001;
		13'b0110101001000: colour_data = 24'b011010101110001101011001;
		13'b0110101001001: colour_data = 24'b011010101110001101011001;
		13'b0110101001010: colour_data = 24'b001000011000111000100001;
		13'b0110101001011: colour_data = 24'b001000011000111000100001;
		13'b0110101001100: colour_data = 24'b000110000110110100011000;
		13'b0110101001101: colour_data = 24'b000110000110110100011000;
		13'b0110101001110: colour_data = 24'b000110000110110100011000;
		13'b0110101001111: colour_data = 24'b000110000110110100011000;
		13'b0110101010000: colour_data = 24'b000110000110110100011000;
		13'b0110101010001: colour_data = 24'b011010101110001101011001;
		13'b0110101010010: colour_data = 24'b011010101110001101011001;
		13'b0110101010011: colour_data = 24'b000110000110110100011000;
		13'b0110101010100: colour_data = 24'b001000011000111000100001;
		13'b0110101010101: colour_data = 24'b001000011000111000100001;
		13'b0110101010110: colour_data = 24'b000110000101000100011000;
		13'b0110101010111: colour_data = 24'b001010101100010100011000;
		13'b0110101011000: colour_data = 24'b000110000110110100011000;
		13'b0110101011001: colour_data = 24'b000110000110110100011000;
		13'b0110101011010: colour_data = 24'b011010101110001101011001;
		13'b0110101011011: colour_data = 24'b011010101110001101011001;
		13'b0110101011100: colour_data = 24'b011010101110001101011001;
		13'b0110101011101: colour_data = 24'b001000011000111000100001;
		13'b0110101011110: colour_data = 24'b001000011000111000100001;
		13'b0110101011111: colour_data = 24'b000110000110110100011000;
		13'b0110101100000: colour_data = 24'b000110000110110100011000;
		13'b0110101100001: colour_data = 24'b000110000110110100011000;
		13'b0110101100010: colour_data = 24'b000110000110110100011000;
		13'b0110101100011: colour_data = 24'b000110000110110100011000;
		13'b0110101100100: colour_data = 24'b011010101110001101011001;
		13'b0110101100101: colour_data = 24'b011010101110001101011001;
		13'b0110101100110: colour_data = 24'b000110000110110100011000;
		13'b0110101100111: colour_data = 24'b001000011000111000100001;
		13'b0110101101000: colour_data = 24'b001000011000111000100001;
		13'b0110101101001: colour_data = 24'b000110000101000100011000;
		13'b0110101101010: colour_data = 24'b001010101100010100011000;
		13'b0110101101011: colour_data = 24'b000110000110110100011000;
		13'b0110101101100: colour_data = 24'b000110000110110100011000;
		13'b0110101101101: colour_data = 24'b011010101110001101011001;
		13'b0110101101110: colour_data = 24'b011010101110001101011001;
		13'b0110101101111: colour_data = 24'b011010101110001101011001;
		13'b0110101110000: colour_data = 24'b001000011000111000100001;
		13'b0110101110001: colour_data = 24'b001000011000111000100001;
		13'b0110101110010: colour_data = 24'b000110000110110100011000;
		13'b0110101110011: colour_data = 24'b000110000110110100011000;
		13'b0110101110100: colour_data = 24'b000110000110110100011000;
		13'b0110101110101: colour_data = 24'b000110000110110100011000;
		13'b0110101110110: colour_data = 24'b000110000110110100011000;
		13'b0110101110111: colour_data = 24'b000110000101000100011000;
		13'b0110101111000: colour_data = 24'b000110000110110100011000;
		13'b0110101111001: colour_data = 24'b000110000110110100011000;
		13'b0110101111010: colour_data = 24'b000110000110110100011000;
		13'b0110101111011: colour_data = 24'b011010101110001101011001;
		13'b0110101111100: colour_data = 24'b011010101110001101011001;
		13'b0110101111101: colour_data = 24'b011010101110001101011001;
		13'b0110101111110: colour_data = 24'b001000011000111000100001;
		13'b0110101111111: colour_data = 24'b001000011000111000100001;
		13'b0110110000000: colour_data = 24'b000110000110110100011000;
		13'b0110110000001: colour_data = 24'b000110000110110100011000;
		13'b0110110000010: colour_data = 24'b001010101100010100011000;
		13'b0110110000011: colour_data = 24'b000110000110110100011000;
		13'b0110110000100: colour_data = 24'b000110000110110100011000;
		13'b0110110000101: colour_data = 24'b011010101110001101011001;
		13'b0110110000110: colour_data = 24'b011010101110001101011001;
		13'b0110110000111: colour_data = 24'b000110000110110100011000;
		13'b0110110001000: colour_data = 24'b111111110000000010010110;
		13'b0110110001001: colour_data = 24'b111111110000000010010110;

		13'b0111000000000: colour_data = 24'b111111110000000010010110;
		13'b0111000000001: colour_data = 24'b111111110000000010010110;
		13'b0111000000010: colour_data = 24'b111111110000000010010110;
		13'b0111000000011: colour_data = 24'b000110000110110100011000;
		13'b0111000000100: colour_data = 24'b000110000110110100011000;
		13'b0111000000101: colour_data = 24'b011010101110001101011001;
		13'b0111000000110: colour_data = 24'b011010101110001101011001;
		13'b0111000000111: colour_data = 24'b000110000110110100011000;
		13'b0111000001000: colour_data = 24'b001000011000111000100001;
		13'b0111000001001: colour_data = 24'b001000011000111000100001;
		13'b0111000001010: colour_data = 24'b000110000101000100011000;
		13'b0111000001011: colour_data = 24'b000110000110110100011000;
		13'b0111000001100: colour_data = 24'b000110000110110100011000;
		13'b0111000001101: colour_data = 24'b000110000110110100011000;
		13'b0111000001110: colour_data = 24'b000110000110110100011000;
		13'b0111000001111: colour_data = 24'b011010101110001101011001;
		13'b0111000010000: colour_data = 24'b001010101100010100011000;
		13'b0111000010001: colour_data = 24'b001000011000111000100001;
		13'b0111000010010: colour_data = 24'b001000011000111000100001;
		13'b0111000010011: colour_data = 24'b011010101110001101011001;
		13'b0111000010100: colour_data = 24'b011010101110001101011001;
		13'b0111000010101: colour_data = 24'b001010101100010100011000;
		13'b0111000010110: colour_data = 24'b001000011000111000100001;
		13'b0111000010111: colour_data = 24'b001000011000111000100001;
		13'b0111000011000: colour_data = 24'b000110000110110100011000;
		13'b0111000011001: colour_data = 24'b000110000110110100011000;
		13'b0111000011010: colour_data = 24'b000110000110110100011000;
		13'b0111000011011: colour_data = 24'b000110000110110100011000;
		13'b0111000011100: colour_data = 24'b000110000110110100011000;
		13'b0111000011101: colour_data = 24'b011010101110001101011001;
		13'b0111000011110: colour_data = 24'b011010101110001101011001;
		13'b0111000011111: colour_data = 24'b000110000110110100011000;
		13'b0111000100000: colour_data = 24'b001000011000111000100001;
		13'b0111000100001: colour_data = 24'b000110000110110100011000;
		13'b0111000100010: colour_data = 24'b000110000101000100011000;
		13'b0111000100011: colour_data = 24'b000110000101000100011000;
		13'b0111000100100: colour_data = 24'b000110000110110100011000;
		13'b0111000100101: colour_data = 24'b000110000110110100011000;
		13'b0111000100110: colour_data = 24'b011010101110001101011001;
		13'b0111000100111: colour_data = 24'b011010101110001101011001;
		13'b0111000101000: colour_data = 24'b001010101100010100011000;
		13'b0111000101001: colour_data = 24'b001000011000111000100001;
		13'b0111000101010: colour_data = 24'b001000011000111000100001;
		13'b0111000101011: colour_data = 24'b000110000110110100011000;
		13'b0111000101100: colour_data = 24'b000110000110110100011000;
		13'b0111000101101: colour_data = 24'b000110000110110100011000;
		13'b0111000101110: colour_data = 24'b000110000110110100011000;
		13'b0111000101111: colour_data = 24'b000110000110110100011000;
		13'b0111000110000: colour_data = 24'b011010101110001101011001;
		13'b0111000110001: colour_data = 24'b001010101100010100011000;
		13'b0111000110010: colour_data = 24'b000110000110110100011000;
		13'b0111000110011: colour_data = 24'b001000011000111000100001;
		13'b0111000110100: colour_data = 24'b000110000110110100011000;
		13'b0111000110101: colour_data = 24'b000110000101000100011000;
		13'b0111000110110: colour_data = 24'b000110000101000100011000;
		13'b0111000110111: colour_data = 24'b000110000110110100011000;
		13'b0111000111000: colour_data = 24'b000110000110110100011000;
		13'b0111000111001: colour_data = 24'b011010101110001101011001;
		13'b0111000111010: colour_data = 24'b011010101110001101011001;
		13'b0111000111011: colour_data = 24'b001010101100010100011000;
		13'b0111000111100: colour_data = 24'b001000011000111000100001;
		13'b0111000111101: colour_data = 24'b001000011000111000100001;
		13'b0111000111110: colour_data = 24'b000110000101000100011000;
		13'b0111000111111: colour_data = 24'b000110000110110100011000;
		13'b0111001000000: colour_data = 24'b000110000110110100011000;
		13'b0111001000001: colour_data = 24'b000110000110110100011000;
		13'b0111001000010: colour_data = 24'b000110000110110100011000;
		13'b0111001000011: colour_data = 24'b011010101110001101011001;
		13'b0111001000100: colour_data = 24'b001010101100010100011000;
		13'b0111001000101: colour_data = 24'b000110000110110100011000;
		13'b0111001000110: colour_data = 24'b001000011000111000100001;
		13'b0111001000111: colour_data = 24'b011010101110001101011001;
		13'b0111001001000: colour_data = 24'b011010101110001101011001;
		13'b0111001001001: colour_data = 24'b001010101100010100011000;
		13'b0111001001010: colour_data = 24'b001000011000111000100001;
		13'b0111001001011: colour_data = 24'b001000011000111000100001;
		13'b0111001001100: colour_data = 24'b000110000110110100011000;
		13'b0111001001101: colour_data = 24'b000110000110110100011000;
		13'b0111001001110: colour_data = 24'b000110000110110100011000;
		13'b0111001001111: colour_data = 24'b000110000110110100011000;
		13'b0111001010000: colour_data = 24'b000110000110110100011000;
		13'b0111001010001: colour_data = 24'b011010101110001101011001;
		13'b0111001010010: colour_data = 24'b011010101110001101011001;
		13'b0111001010011: colour_data = 24'b000110000110110100011000;
		13'b0111001010100: colour_data = 24'b001000011000111000100001;
		13'b0111001010101: colour_data = 24'b001000011000111000100001;
		13'b0111001010110: colour_data = 24'b000110000101000100011000;
		13'b0111001010111: colour_data = 24'b000110000101000100011000;
		13'b0111001011000: colour_data = 24'b000110000110110100011000;
		13'b0111001011001: colour_data = 24'b000110000110110100011000;
		13'b0111001011010: colour_data = 24'b011010101110001101011001;
		13'b0111001011011: colour_data = 24'b011010101110001101011001;
		13'b0111001011100: colour_data = 24'b001010101100010100011000;
		13'b0111001011101: colour_data = 24'b001000011000111000100001;
		13'b0111001011110: colour_data = 24'b001000011000111000100001;
		13'b0111001011111: colour_data = 24'b000110000110110100011000;
		13'b0111001100000: colour_data = 24'b000110000110110100011000;
		13'b0111001100001: colour_data = 24'b000110000110110100011000;
		13'b0111001100010: colour_data = 24'b000110000110110100011000;
		13'b0111001100011: colour_data = 24'b000110000110110100011000;
		13'b0111001100100: colour_data = 24'b011010101110001101011001;
		13'b0111001100101: colour_data = 24'b011010101110001101011001;
		13'b0111001100110: colour_data = 24'b000110000110110100011000;
		13'b0111001100111: colour_data = 24'b001000011000111000100001;
		13'b0111001101000: colour_data = 24'b001000011000111000100001;
		13'b0111001101001: colour_data = 24'b000110000101000100011000;
		13'b0111001101010: colour_data = 24'b000110000101000100011000;
		13'b0111001101011: colour_data = 24'b000110000110110100011000;
		13'b0111001101100: colour_data = 24'b000110000110110100011000;
		13'b0111001101101: colour_data = 24'b011010101110001101011001;
		13'b0111001101110: colour_data = 24'b011010101110001101011001;
		13'b0111001101111: colour_data = 24'b001010101100010100011000;
		13'b0111001110000: colour_data = 24'b001000011000111000100001;
		13'b0111001110001: colour_data = 24'b001000011000111000100001;
		13'b0111001110010: colour_data = 24'b000110000110110100011000;
		13'b0111001110011: colour_data = 24'b000110000110110100011000;
		13'b0111001110100: colour_data = 24'b000110000110110100011000;
		13'b0111001110101: colour_data = 24'b000110000110110100011000;
		13'b0111001110110: colour_data = 24'b000110000110110100011000;
		13'b0111001110111: colour_data = 24'b000110000101000100011000;
		13'b0111001111000: colour_data = 24'b000110000110110100011000;
		13'b0111001111001: colour_data = 24'b000110000110110100011000;
		13'b0111001111010: colour_data = 24'b000110000110110100011000;
		13'b0111001111011: colour_data = 24'b011010101110001101011001;
		13'b0111001111100: colour_data = 24'b011010101110001101011001;
		13'b0111001111101: colour_data = 24'b001010101100010100011000;
		13'b0111001111110: colour_data = 24'b001000011000111000100001;
		13'b0111001111111: colour_data = 24'b001000011000111000100001;
		13'b0111010000000: colour_data = 24'b000110000110110100011000;
		13'b0111010000001: colour_data = 24'b000110000110110100011000;
		13'b0111010000010: colour_data = 24'b000110000101000100011000;
		13'b0111010000011: colour_data = 24'b000110000110110100011000;
		13'b0111010000100: colour_data = 24'b000110000110110100011000;
		13'b0111010000101: colour_data = 24'b011010101110001101011001;
		13'b0111010000110: colour_data = 24'b011010101110001101011001;
		13'b0111010000111: colour_data = 24'b111111110000000010010110;
		13'b0111010001000: colour_data = 24'b111111110000000010010110;
		13'b0111010001001: colour_data = 24'b111111110000000010010110;

		13'b0111100000000: colour_data = 24'b111111110000000010010110;
		13'b0111100000001: colour_data = 24'b111111110000000010010110;
		13'b0111100000010: colour_data = 24'b111111110000000010010110;
		13'b0111100000011: colour_data = 24'b000110000110110100011000;
		13'b0111100000100: colour_data = 24'b000110000110110100011000;
		13'b0111100000101: colour_data = 24'b011010101110001101011001;
		13'b0111100000110: colour_data = 24'b011010101110001101011001;
		13'b0111100000111: colour_data = 24'b000110000110110100011000;
		13'b0111100001000: colour_data = 24'b001000011000111000100001;
		13'b0111100001001: colour_data = 24'b001000011000111000100001;
		13'b0111100001010: colour_data = 24'b000110000101000100011000;
		13'b0111100001011: colour_data = 24'b000110000110110100011000;
		13'b0111100001100: colour_data = 24'b000110000110110100011000;
		13'b0111100001101: colour_data = 24'b000110000110110100011000;
		13'b0111100001110: colour_data = 24'b000110000110110100011000;
		13'b0111100001111: colour_data = 24'b001010101100010100011000;
		13'b0111100010000: colour_data = 24'b001010101100010100011000;
		13'b0111100010001: colour_data = 24'b001000011000111000100001;
		13'b0111100010010: colour_data = 24'b001000011000111000100001;
		13'b0111100010011: colour_data = 24'b011010101110001101011001;
		13'b0111100010100: colour_data = 24'b011010101110001101011001;
		13'b0111100010101: colour_data = 24'b001010101100010100011000;
		13'b0111100010110: colour_data = 24'b001000011000111000100001;
		13'b0111100010111: colour_data = 24'b001000011000111000100001;
		13'b0111100011000: colour_data = 24'b000110000110110100011000;
		13'b0111100011001: colour_data = 24'b000110000110110100011000;
		13'b0111100011010: colour_data = 24'b000110000110110100011000;
		13'b0111100011011: colour_data = 24'b000110000110110100011000;
		13'b0111100011100: colour_data = 24'b000110000110110100011000;
		13'b0111100011101: colour_data = 24'b001010101100010100011000;
		13'b0111100011110: colour_data = 24'b011010101110001101011001;
		13'b0111100011111: colour_data = 24'b000110000110110100011000;
		13'b0111100100000: colour_data = 24'b001000011000111000100001;
		13'b0111100100001: colour_data = 24'b000110000110110100011000;
		13'b0111100100010: colour_data = 24'b000110000101000100011000;
		13'b0111100100011: colour_data = 24'b000110000101000100011000;
		13'b0111100100100: colour_data = 24'b000110000110110100011000;
		13'b0111100100101: colour_data = 24'b000110000110110100011000;
		13'b0111100100110: colour_data = 24'b011010101110001101011001;
		13'b0111100100111: colour_data = 24'b011010101110001101011001;
		13'b0111100101000: colour_data = 24'b001010101100010100011000;
		13'b0111100101001: colour_data = 24'b001000011000111000100001;
		13'b0111100101010: colour_data = 24'b001000011000111000100001;
		13'b0111100101011: colour_data = 24'b000110000110110100011000;
		13'b0111100101100: colour_data = 24'b000110000110110100011000;
		13'b0111100101101: colour_data = 24'b000110000110110100011000;
		13'b0111100101110: colour_data = 24'b000110000110110100011000;
		13'b0111100101111: colour_data = 24'b000110000110110100011000;
		13'b0111100110000: colour_data = 24'b001010101100010100011000;
		13'b0111100110001: colour_data = 24'b001010101100010100011000;
		13'b0111100110010: colour_data = 24'b000110000110110100011000;
		13'b0111100110011: colour_data = 24'b001000011000111000100001;
		13'b0111100110100: colour_data = 24'b000110000110110100011000;
		13'b0111100110101: colour_data = 24'b000110000101000100011000;
		13'b0111100110110: colour_data = 24'b000110000101000100011000;
		13'b0111100110111: colour_data = 24'b000110000110110100011000;
		13'b0111100111000: colour_data = 24'b000110000110110100011000;
		13'b0111100111001: colour_data = 24'b011010101110001101011001;
		13'b0111100111010: colour_data = 24'b011010101110001101011001;
		13'b0111100111011: colour_data = 24'b001010101100010100011000;
		13'b0111100111100: colour_data = 24'b001000011000111000100001;
		13'b0111100111101: colour_data = 24'b001000011000111000100001;
		13'b0111100111110: colour_data = 24'b000110000101000100011000;
		13'b0111100111111: colour_data = 24'b000110000110110100011000;
		13'b0111101000000: colour_data = 24'b000110000110110100011000;
		13'b0111101000001: colour_data = 24'b000110000110110100011000;
		13'b0111101000010: colour_data = 24'b000110000110110100011000;
		13'b0111101000011: colour_data = 24'b001010101100010100011000;
		13'b0111101000100: colour_data = 24'b001010101100010100011000;
		13'b0111101000101: colour_data = 24'b000110000110110100011000;
		13'b0111101000110: colour_data = 24'b001000011000111000100001;
		13'b0111101000111: colour_data = 24'b011010101110001101011001;
		13'b0111101001000: colour_data = 24'b001010101100010100011000;
		13'b0111101001001: colour_data = 24'b001010101100010100011000;
		13'b0111101001010: colour_data = 24'b001000011000111000100001;
		13'b0111101001011: colour_data = 24'b001000011000111000100001;
		13'b0111101001100: colour_data = 24'b000110000110110100011000;
		13'b0111101001101: colour_data = 24'b000110000110110100011000;
		13'b0111101001110: colour_data = 24'b000110000110110100011000;
		13'b0111101001111: colour_data = 24'b000110000110110100011000;
		13'b0111101010000: colour_data = 24'b000110000110110100011000;
		13'b0111101010001: colour_data = 24'b001010101100010100011000;
		13'b0111101010010: colour_data = 24'b011010101110001101011001;
		13'b0111101010011: colour_data = 24'b000110000110110100011000;
		13'b0111101010100: colour_data = 24'b001000011000111000100001;
		13'b0111101010101: colour_data = 24'b001000011000111000100001;
		13'b0111101010110: colour_data = 24'b000110000101000100011000;
		13'b0111101010111: colour_data = 24'b000110000101000100011000;
		13'b0111101011000: colour_data = 24'b000110000110110100011000;
		13'b0111101011001: colour_data = 24'b000110000110110100011000;
		13'b0111101011010: colour_data = 24'b011010101110001101011001;
		13'b0111101011011: colour_data = 24'b001010101100010100011000;
		13'b0111101011100: colour_data = 24'b001010101100010100011000;
		13'b0111101011101: colour_data = 24'b001000011000111000100001;
		13'b0111101011110: colour_data = 24'b001000011000111000100001;
		13'b0111101011111: colour_data = 24'b000110000110110100011000;
		13'b0111101100000: colour_data = 24'b000110000110110100011000;
		13'b0111101100001: colour_data = 24'b000110000110110100011000;
		13'b0111101100010: colour_data = 24'b000110000110110100011000;
		13'b0111101100011: colour_data = 24'b000110000110110100011000;
		13'b0111101100100: colour_data = 24'b001010101100010100011000;
		13'b0111101100101: colour_data = 24'b011010101110001101011001;
		13'b0111101100110: colour_data = 24'b000110000110110100011000;
		13'b0111101100111: colour_data = 24'b001000011000111000100001;
		13'b0111101101000: colour_data = 24'b001000011000111000100001;
		13'b0111101101001: colour_data = 24'b000110000101000100011000;
		13'b0111101101010: colour_data = 24'b000110000101000100011000;
		13'b0111101101011: colour_data = 24'b000110000110110100011000;
		13'b0111101101100: colour_data = 24'b000110000110110100011000;
		13'b0111101101101: colour_data = 24'b011010101110001101011001;
		13'b0111101101110: colour_data = 24'b011010101110001101011001;
		13'b0111101101111: colour_data = 24'b001010101100010100011000;
		13'b0111101110000: colour_data = 24'b001000011000111000100001;
		13'b0111101110001: colour_data = 24'b001000011000111000100001;
		13'b0111101110010: colour_data = 24'b000110000110110100011000;
		13'b0111101110011: colour_data = 24'b000110000110110100011000;
		13'b0111101110100: colour_data = 24'b000110000110110100011000;
		13'b0111101110101: colour_data = 24'b000110000110110100011000;
		13'b0111101110110: colour_data = 24'b000110000110110100011000;
		13'b0111101110111: colour_data = 24'b000110000101000100011000;
		13'b0111101111000: colour_data = 24'b000110000110110100011000;
		13'b0111101111001: colour_data = 24'b000110000110110100011000;
		13'b0111101111010: colour_data = 24'b000110000110110100011000;
		13'b0111101111011: colour_data = 24'b011010101110001101011001;
		13'b0111101111100: colour_data = 24'b001010101100010100011000;
		13'b0111101111101: colour_data = 24'b001010101100010100011000;
		13'b0111101111110: colour_data = 24'b001000011000111000100001;
		13'b0111101111111: colour_data = 24'b001000011000111000100001;
		13'b0111110000000: colour_data = 24'b000110000110110100011000;
		13'b0111110000001: colour_data = 24'b000110000110110100011000;
		13'b0111110000010: colour_data = 24'b000110000101000100011000;
		13'b0111110000011: colour_data = 24'b000110000110110100011000;
		13'b0111110000100: colour_data = 24'b000110000110110100011000;
		13'b0111110000101: colour_data = 24'b011010101110001101011001;
		13'b0111110000110: colour_data = 24'b011010101110001101011001;
		13'b0111110000111: colour_data = 24'b111111110000000010010110;
		13'b0111110001000: colour_data = 24'b111111110000000010010110;
		13'b0111110001001: colour_data = 24'b111111110000000010010110;

		13'b1000000000000: colour_data = 24'b111111110000000010010110;
		13'b1000000000001: colour_data = 24'b111111110000000010010110;
		13'b1000000000010: colour_data = 24'b111111110000000010010110;
		13'b1000000000011: colour_data = 24'b000110000110110100011000;
		13'b1000000000100: colour_data = 24'b000110000110110100011000;
		13'b1000000000101: colour_data = 24'b011010101110001101011001;
		13'b1000000000110: colour_data = 24'b001010101100010100011000;
		13'b1000000000111: colour_data = 24'b111111110000000010010110;
		13'b1000000001000: colour_data = 24'b000110000110110100011000;
		13'b1000000001001: colour_data = 24'b001000011000111000100001;
		13'b1000000001010: colour_data = 24'b000110000101000100011000;
		13'b1000000001011: colour_data = 24'b000110000101000100011000;
		13'b1000000001100: colour_data = 24'b111111110000000010010110;
		13'b1000000001101: colour_data = 24'b000110000110110100011000;
		13'b1000000001110: colour_data = 24'b000110000110110100011000;
		13'b1000000001111: colour_data = 24'b001010101100010100011000;
		13'b1000000010000: colour_data = 24'b111111110000000010010110;
		13'b1000000010001: colour_data = 24'b000110000110110100011000;
		13'b1000000010010: colour_data = 24'b001000011000111000100001;
		13'b1000000010011: colour_data = 24'b011010101110001101011001;
		13'b1000000010100: colour_data = 24'b001010101100010100011000;
		13'b1000000010101: colour_data = 24'b111111110000000010010110;
		13'b1000000010110: colour_data = 24'b000110000110110100011000;
		13'b1000000010111: colour_data = 24'b001000011000111000100001;
		13'b1000000011000: colour_data = 24'b000110000110110100011000;
		13'b1000000011001: colour_data = 24'b000110000101000100011000;
		13'b1000000011010: colour_data = 24'b111111110000000010010110;
		13'b1000000011011: colour_data = 24'b000110000110110100011000;
		13'b1000000011100: colour_data = 24'b000110000110110100011000;
		13'b1000000011101: colour_data = 24'b001010101100010100011000;
		13'b1000000011110: colour_data = 24'b001010101100010100011000;
		13'b1000000011111: colour_data = 24'b111111110000000010010110;
		13'b1000000100000: colour_data = 24'b001000011000111000100001;
		13'b1000000100001: colour_data = 24'b000110000110110100011000;
		13'b1000000100010: colour_data = 24'b000110000101000100011000;
		13'b1000000100011: colour_data = 24'b111111110000000010010110;
		13'b1000000100100: colour_data = 24'b000110000110110100011000;
		13'b1000000100101: colour_data = 24'b000110000110110100011000;
		13'b1000000100110: colour_data = 24'b011010101110001101011001;
		13'b1000000100111: colour_data = 24'b001010101100010100011000;
		13'b1000000101000: colour_data = 24'b111111110000000010010110;
		13'b1000000101001: colour_data = 24'b000110000110110100011000;
		13'b1000000101010: colour_data = 24'b001000011000111000100001;
		13'b1000000101011: colour_data = 24'b000110000110110100011000;
		13'b1000000101100: colour_data = 24'b000110000101000100011000;
		13'b1000000101101: colour_data = 24'b111111110000000010010110;
		13'b1000000101110: colour_data = 24'b000110000110110100011000;
		13'b1000000101111: colour_data = 24'b000110000110110100011000;
		13'b1000000110000: colour_data = 24'b001010101100010100011000;
		13'b1000000110001: colour_data = 24'b111111110000000010010110;
		13'b1000000110010: colour_data = 24'b111111110000000010010110;
		13'b1000000110011: colour_data = 24'b001000011000111000100001;
		13'b1000000110100: colour_data = 24'b000110000110110100011000;
		13'b1000000110101: colour_data = 24'b000110000101000100011000;
		13'b1000000110110: colour_data = 24'b111111110000000010010110;
		13'b1000000110111: colour_data = 24'b000110000110110100011000;
		13'b1000000111000: colour_data = 24'b000110000110110100011000;
		13'b1000000111001: colour_data = 24'b011010101110001101011001;
		13'b1000000111010: colour_data = 24'b001010101100010100011000;
		13'b1000000111011: colour_data = 24'b111111110000000010010110;
		13'b1000000111100: colour_data = 24'b000110000110110100011000;
		13'b1000000111101: colour_data = 24'b001000011000111000100001;
		13'b1000000111110: colour_data = 24'b000110000101000100011000;
		13'b1000000111111: colour_data = 24'b000110000101000100011000;
		13'b1000001000000: colour_data = 24'b111111110000000010010110;
		13'b1000001000001: colour_data = 24'b000110000110110100011000;
		13'b1000001000010: colour_data = 24'b000110000110110100011000;
		13'b1000001000011: colour_data = 24'b001010101100010100011000;
		13'b1000001000100: colour_data = 24'b111111110000000010010110;
		13'b1000001000101: colour_data = 24'b111111110000000010010110;
		13'b1000001000110: colour_data = 24'b001000011000111000100001;
		13'b1000001000111: colour_data = 24'b011010101110001101011001;
		13'b1000001001000: colour_data = 24'b001010101100010100011000;
		13'b1000001001001: colour_data = 24'b111111110000000010010110;
		13'b1000001001010: colour_data = 24'b000110000110110100011000;
		13'b1000001001011: colour_data = 24'b001000011000111000100001;
		13'b1000001001100: colour_data = 24'b000110000110110100011000;
		13'b1000001001101: colour_data = 24'b000110000101000100011000;
		13'b1000001001110: colour_data = 24'b111111110000000010010110;
		13'b1000001001111: colour_data = 24'b000110000110110100011000;
		13'b1000001010000: colour_data = 24'b000110000110110100011000;
		13'b1000001010001: colour_data = 24'b001010101100010100011000;
		13'b1000001010010: colour_data = 24'b001010101100010100011000;
		13'b1000001010011: colour_data = 24'b111111110000000010010110;
		13'b1000001010100: colour_data = 24'b001000011000111000100001;
		13'b1000001010101: colour_data = 24'b001000011000111000100001;
		13'b1000001010110: colour_data = 24'b000110000101000100011000;
		13'b1000001010111: colour_data = 24'b111111110000000010010110;
		13'b1000001011000: colour_data = 24'b111111110000000010010110;
		13'b1000001011001: colour_data = 24'b000110000110110100011000;
		13'b1000001011010: colour_data = 24'b011010101110001101011001;
		13'b1000001011011: colour_data = 24'b001010101100010100011000;
		13'b1000001011100: colour_data = 24'b111111110000000010010110;
		13'b1000001011101: colour_data = 24'b000110000110110100011000;
		13'b1000001011110: colour_data = 24'b001000011000111000100001;
		13'b1000001011111: colour_data = 24'b000110000110110100011000;
		13'b1000001100000: colour_data = 24'b000110000101000100011000;
		13'b1000001100001: colour_data = 24'b111111110000000010010110;
		13'b1000001100010: colour_data = 24'b000110000110110100011000;
		13'b1000001100011: colour_data = 24'b000110000110110100011000;
		13'b1000001100100: colour_data = 24'b001010101100010100011000;
		13'b1000001100101: colour_data = 24'b001010101100010100011000;
		13'b1000001100110: colour_data = 24'b111111110000000010010110;
		13'b1000001100111: colour_data = 24'b001000011000111000100001;
		13'b1000001101000: colour_data = 24'b001000011000111000100001;
		13'b1000001101001: colour_data = 24'b000110000101000100011000;
		13'b1000001101010: colour_data = 24'b111111110000000010010110;
		13'b1000001101011: colour_data = 24'b000110000110110100011000;
		13'b1000001101100: colour_data = 24'b000110000110110100011000;
		13'b1000001101101: colour_data = 24'b011010101110001101011001;
		13'b1000001101110: colour_data = 24'b001010101100010100011000;
		13'b1000001101111: colour_data = 24'b111111110000000010010110;
		13'b1000001110000: colour_data = 24'b000110000110110100011000;
		13'b1000001110001: colour_data = 24'b001000011000111000100001;
		13'b1000001110010: colour_data = 24'b000110000110110100011000;
		13'b1000001110011: colour_data = 24'b000110000101000100011000;
		13'b1000001110100: colour_data = 24'b111111110000000010010110;
		13'b1000001110101: colour_data = 24'b000110000110110100011000;
		13'b1000001110110: colour_data = 24'b000110000110110100011000;
		13'b1000001110111: colour_data = 24'b000110000101000100011000;
		13'b1000001111000: colour_data = 24'b000110000101000100011000;
		13'b1000001111001: colour_data = 24'b111111110000000010010110;
		13'b1000001111010: colour_data = 24'b000110000110110100011000;
		13'b1000001111011: colour_data = 24'b011010101110001101011001;
		13'b1000001111100: colour_data = 24'b001010101100010100011000;
		13'b1000001111101: colour_data = 24'b111111110000000010010110;
		13'b1000001111110: colour_data = 24'b000110000110110100011000;
		13'b1000001111111: colour_data = 24'b001000011000111000100001;
		13'b1000010000000: colour_data = 24'b000110000110110100011000;
		13'b1000010000001: colour_data = 24'b000110000101000100011000;
		13'b1000010000010: colour_data = 24'b111111110000000010010110;
		13'b1000010000011: colour_data = 24'b000110000110110100011000;
		13'b1000010000100: colour_data = 24'b000110000110110100011000;
		13'b1000010000101: colour_data = 24'b011010101110001101011001;
		13'b1000010000110: colour_data = 24'b001010101100010100011000;
		13'b1000010000111: colour_data = 24'b111111110000000010010110;
		13'b1000010001000: colour_data = 24'b111111110000000010010110;
		13'b1000010001001: colour_data = 24'b111111110000000010010110;

		13'b1000100000000: colour_data = 24'b111111110000000010010110;
		13'b1000100000001: colour_data = 24'b111111110000000010010110;
		13'b1000100000010: colour_data = 24'b111111110000000010010110;
		13'b1000100000011: colour_data = 24'b111111110000000010010110;
		13'b1000100000100: colour_data = 24'b000110000110110100011000;
		13'b1000100000101: colour_data = 24'b011010101110001101011001;
		13'b1000100000110: colour_data = 24'b111111110000000010010110;
		13'b1000100000111: colour_data = 24'b111111110000000010010110;
		13'b1000100001000: colour_data = 24'b111111110000000010010110;
		13'b1000100001001: colour_data = 24'b001000011000111000100001;
		13'b1000100001010: colour_data = 24'b000110000101000100011000;
		13'b1000100001011: colour_data = 24'b111111110000000010010110;
		13'b1000100001100: colour_data = 24'b111111110000000010010110;
		13'b1000100001101: colour_data = 24'b000110000110110100011000;
		13'b1000100001110: colour_data = 24'b000110000110110100011000;
		13'b1000100001111: colour_data = 24'b000110000101000100011000;
		13'b1000100010000: colour_data = 24'b111111110000000010010110;
		13'b1000100010001: colour_data = 24'b111111110000000010010110;
		13'b1000100010010: colour_data = 24'b000110000110110100011000;
		13'b1000100010011: colour_data = 24'b011010101110001101011001;
		13'b1000100010100: colour_data = 24'b111111110000000010010110;
		13'b1000100010101: colour_data = 24'b111111110000000010010110;
		13'b1000100010110: colour_data = 24'b111111110000000010010110;
		13'b1000100010111: colour_data = 24'b001000011000111000100001;
		13'b1000100011000: colour_data = 24'b000110000101000100011000;
		13'b1000100011001: colour_data = 24'b111111110000000010010110;
		13'b1000100011010: colour_data = 24'b111111110000000010010110;
		13'b1000100011011: colour_data = 24'b111111110000000010010110;
		13'b1000100011100: colour_data = 24'b000110000110110100011000;
		13'b1000100011101: colour_data = 24'b001010101100010100011000;
		13'b1000100011110: colour_data = 24'b111111110000000010010110;
		13'b1000100011111: colour_data = 24'b111111110000000010010110;
		13'b1000100100000: colour_data = 24'b000110000110110100011000;
		13'b1000100100001: colour_data = 24'b000110000101000100011000;
		13'b1000100100010: colour_data = 24'b000110000101000100011000;
		13'b1000100100011: colour_data = 24'b111111110000000010010110;
		13'b1000100100100: colour_data = 24'b111111110000000010010110;
		13'b1000100100101: colour_data = 24'b000110000110110100011000;
		13'b1000100100110: colour_data = 24'b011010101110001101011001;
		13'b1000100100111: colour_data = 24'b111111110000000010010110;
		13'b1000100101000: colour_data = 24'b111111110000000010010110;
		13'b1000100101001: colour_data = 24'b111111110000000010010110;
		13'b1000100101010: colour_data = 24'b001000011000111000100001;
		13'b1000100101011: colour_data = 24'b000110000101000100011000;
		13'b1000100101100: colour_data = 24'b111111110000000010010110;
		13'b1000100101101: colour_data = 24'b111111110000000010010110;
		13'b1000100101110: colour_data = 24'b111111110000000010010110;
		13'b1000100101111: colour_data = 24'b000110000110110100011000;
		13'b1000100110000: colour_data = 24'b001010101100010100011000;
		13'b1000100110001: colour_data = 24'b111111110000000010010110;
		13'b1000100110010: colour_data = 24'b111111110000000010010110;
		13'b1000100110011: colour_data = 24'b000110000110110100011000;
		13'b1000100110100: colour_data = 24'b000110000101000100011000;
		13'b1000100110101: colour_data = 24'b000110000101000100011000;
		13'b1000100110110: colour_data = 24'b111111110000000010010110;
		13'b1000100110111: colour_data = 24'b111111110000000010010110;
		13'b1000100111000: colour_data = 24'b000110000110110100011000;
		13'b1000100111001: colour_data = 24'b011010101110001101011001;
		13'b1000100111010: colour_data = 24'b111111110000000010010110;
		13'b1000100111011: colour_data = 24'b111111110000000010010110;
		13'b1000100111100: colour_data = 24'b111111110000000010010110;
		13'b1000100111101: colour_data = 24'b001000011000111000100001;
		13'b1000100111110: colour_data = 24'b000110000101000100011000;
		13'b1000100111111: colour_data = 24'b111111110000000010010110;
		13'b1000101000000: colour_data = 24'b111111110000000010010110;
		13'b1000101000001: colour_data = 24'b000110000110110100011000;
		13'b1000101000010: colour_data = 24'b000110000110110100011000;
		13'b1000101000011: colour_data = 24'b000110000101000100011000;
		13'b1000101000100: colour_data = 24'b111111110000000010010110;
		13'b1000101000101: colour_data = 24'b111111110000000010010110;
		13'b1000101000110: colour_data = 24'b000110000110110100011000;
		13'b1000101000111: colour_data = 24'b011010101110001101011001;
		13'b1000101001000: colour_data = 24'b001010101100010100011000;
		13'b1000101001001: colour_data = 24'b111111110000000010010110;
		13'b1000101001010: colour_data = 24'b111111110000000010010110;
		13'b1000101001011: colour_data = 24'b000110000110110100011000;
		13'b1000101001100: colour_data = 24'b000110000101000100011000;
		13'b1000101001101: colour_data = 24'b111111110000000010010110;
		13'b1000101001110: colour_data = 24'b111111110000000010010110;
		13'b1000101001111: colour_data = 24'b111111110000000010010110;
		13'b1000101010000: colour_data = 24'b000110000110110100011000;
		13'b1000101010001: colour_data = 24'b001010101100010100011000;
		13'b1000101010010: colour_data = 24'b111111110000000010010110;
		13'b1000101010011: colour_data = 24'b111111110000000010010110;
		13'b1000101010100: colour_data = 24'b000110000110110100011000;
		13'b1000101010101: colour_data = 24'b001000011000111000100001;
		13'b1000101010110: colour_data = 24'b000110000101000100011000;
		13'b1000101010111: colour_data = 24'b111111110000000010010110;
		13'b1000101011000: colour_data = 24'b111111110000000010010110;
		13'b1000101011001: colour_data = 24'b000110000110110100011000;
		13'b1000101011010: colour_data = 24'b011010101110001101011001;
		13'b1000101011011: colour_data = 24'b001010101100010100011000;
		13'b1000101011100: colour_data = 24'b111111110000000010010110;
		13'b1000101011101: colour_data = 24'b111111110000000010010110;
		13'b1000101011110: colour_data = 24'b001000011000111000100001;
		13'b1000101011111: colour_data = 24'b000110000101000100011000;
		13'b1000101100000: colour_data = 24'b111111110000000010010110;
		13'b1000101100001: colour_data = 24'b111111110000000010010110;
		13'b1000101100010: colour_data = 24'b111111110000000010010110;
		13'b1000101100011: colour_data = 24'b000110000110110100011000;
		13'b1000101100100: colour_data = 24'b001010101100010100011000;
		13'b1000101100101: colour_data = 24'b111111110000000010010110;
		13'b1000101100110: colour_data = 24'b111111110000000010010110;
		13'b1000101100111: colour_data = 24'b000110000110110100011000;
		13'b1000101101000: colour_data = 24'b001000011000111000100001;
		13'b1000101101001: colour_data = 24'b000110000101000100011000;
		13'b1000101101010: colour_data = 24'b111111110000000010010110;
		13'b1000101101011: colour_data = 24'b111111110000000010010110;
		13'b1000101101100: colour_data = 24'b000110000110110100011000;
		13'b1000101101101: colour_data = 24'b011010101110001101011001;
		13'b1000101101110: colour_data = 24'b111111110000000010010110;
		13'b1000101101111: colour_data = 24'b111111110000000010010110;
		13'b1000101110000: colour_data = 24'b111111110000000010010110;
		13'b1000101110001: colour_data = 24'b001000011000111000100001;
		13'b1000101110010: colour_data = 24'b000110000101000100011000;
		13'b1000101110011: colour_data = 24'b111111110000000010010110;
		13'b1000101110100: colour_data = 24'b111111110000000010010110;
		13'b1000101110101: colour_data = 24'b111111110000000010010110;
		13'b1000101110110: colour_data = 24'b000110000110110100011000;
		13'b1000101110111: colour_data = 24'b000110000101000100011000;
		13'b1000101111000: colour_data = 24'b111111110000000010010110;
		13'b1000101111001: colour_data = 24'b111111110000000010010110;
		13'b1000101111010: colour_data = 24'b000110000110110100011000;
		13'b1000101111011: colour_data = 24'b011010101110001101011001;
		13'b1000101111100: colour_data = 24'b001010101100010100011000;
		13'b1000101111101: colour_data = 24'b111111110000000010010110;
		13'b1000101111110: colour_data = 24'b111111110000000010010110;
		13'b1000101111111: colour_data = 24'b000110000110110100011000;
		13'b1000110000000: colour_data = 24'b000110000101000100011000;
		13'b1000110000001: colour_data = 24'b111111110000000010010110;
		13'b1000110000010: colour_data = 24'b111111110000000010010110;
		13'b1000110000011: colour_data = 24'b111111110000000010010110;
		13'b1000110000100: colour_data = 24'b000110000110110100011000;
		13'b1000110000101: colour_data = 24'b011010101110001101011001;
		13'b1000110000110: colour_data = 24'b111111110000000010010110;
		13'b1000110000111: colour_data = 24'b111111110000000010010110;
		13'b1000110001000: colour_data = 24'b111111110000000010010110;
		13'b1000110001001: colour_data = 24'b111111110000000010010110;

		13'b1001000000000: colour_data = 24'b111111110000000010010110;
		13'b1001000000001: colour_data = 24'b111111110000000010010110;
		13'b1001000000010: colour_data = 24'b111111110000000010010110;
		13'b1001000000011: colour_data = 24'b111111110000000010010110;
		13'b1001000000100: colour_data = 24'b000110000110110100011000;
		13'b1001000000101: colour_data = 24'b001010101100010100011000;
		13'b1001000000110: colour_data = 24'b111111110000000010010110;
		13'b1001000000111: colour_data = 24'b111111110000000010010110;
		13'b1001000001000: colour_data = 24'b111111110000000010010110;
		13'b1001000001001: colour_data = 24'b000110000110110100011000;
		13'b1001000001010: colour_data = 24'b111111110000000010010110;
		13'b1001000001011: colour_data = 24'b111111110000000010010110;
		13'b1001000001100: colour_data = 24'b111111110000000010010110;
		13'b1001000001101: colour_data = 24'b111111110000000010010110;
		13'b1001000001110: colour_data = 24'b000110000110110100011000;
		13'b1001000001111: colour_data = 24'b111111110000000010010110;
		13'b1001000010000: colour_data = 24'b111111110000000010010110;
		13'b1001000010001: colour_data = 24'b111111110000000010010110;
		13'b1001000010010: colour_data = 24'b111111110000000010010110;
		13'b1001000010011: colour_data = 24'b001010101100010100011000;
		13'b1001000010100: colour_data = 24'b111111110000000010010110;
		13'b1001000010101: colour_data = 24'b111111110000000010010110;
		13'b1001000010110: colour_data = 24'b111111110000000010010110;
		13'b1001000010111: colour_data = 24'b000110000110110100011000;
		13'b1001000011000: colour_data = 24'b000110000101000100011000;
		13'b1001000011001: colour_data = 24'b111111110000000010010110;
		13'b1001000011010: colour_data = 24'b111111110000000010010110;
		13'b1001000011011: colour_data = 24'b111111110000000010010110;
		13'b1001000011100: colour_data = 24'b000110000110110100011000;
		13'b1001000011101: colour_data = 24'b111111110000000010010110;
		13'b1001000011110: colour_data = 24'b111111110000000010010110;
		13'b1001000011111: colour_data = 24'b111111110000000010010110;
		13'b1001000100000: colour_data = 24'b111111110000000010010110;
		13'b1001000100001: colour_data = 24'b000110000101000100011000;
		13'b1001000100010: colour_data = 24'b111111110000000010010110;
		13'b1001000100011: colour_data = 24'b111111110000000010010110;
		13'b1001000100100: colour_data = 24'b111111110000000010010110;
		13'b1001000100101: colour_data = 24'b111111110000000010010110;
		13'b1001000100110: colour_data = 24'b001010101100010100011000;
		13'b1001000100111: colour_data = 24'b111111110000000010010110;
		13'b1001000101000: colour_data = 24'b111111110000000010010110;
		13'b1001000101001: colour_data = 24'b111111110000000010010110;
		13'b1001000101010: colour_data = 24'b000110000110110100011000;
		13'b1001000101011: colour_data = 24'b000110000101000100011000;
		13'b1001000101100: colour_data = 24'b111111110000000010010110;
		13'b1001000101101: colour_data = 24'b111111110000000010010110;
		13'b1001000101110: colour_data = 24'b111111110000000010010110;
		13'b1001000101111: colour_data = 24'b000110000110110100011000;
		13'b1001000110000: colour_data = 24'b111111110000000010010110;
		13'b1001000110001: colour_data = 24'b111111110000000010010110;
		13'b1001000110010: colour_data = 24'b111111110000000010010110;
		13'b1001000110011: colour_data = 24'b111111110000000010010110;
		13'b1001000110100: colour_data = 24'b000110000101000100011000;
		13'b1001000110101: colour_data = 24'b111111110000000010010110;
		13'b1001000110110: colour_data = 24'b111111110000000010010110;
		13'b1001000110111: colour_data = 24'b111111110000000010010110;
		13'b1001000111000: colour_data = 24'b111111110000000010010110;
		13'b1001000111001: colour_data = 24'b001010101100010100011000;
		13'b1001000111010: colour_data = 24'b111111110000000010010110;
		13'b1001000111011: colour_data = 24'b111111110000000010010110;
		13'b1001000111100: colour_data = 24'b111111110000000010010110;
		13'b1001000111101: colour_data = 24'b000110000110110100011000;
		13'b1001000111110: colour_data = 24'b111111110000000010010110;
		13'b1001000111111: colour_data = 24'b111111110000000010010110;
		13'b1001001000000: colour_data = 24'b111111110000000010010110;
		13'b1001001000001: colour_data = 24'b111111110000000010010110;
		13'b1001001000010: colour_data = 24'b000110000110110100011000;
		13'b1001001000011: colour_data = 24'b111111110000000010010110;
		13'b1001001000100: colour_data = 24'b111111110000000010010110;
		13'b1001001000101: colour_data = 24'b111111110000000010010110;
		13'b1001001000110: colour_data = 24'b111111110000000010010110;
		13'b1001001000111: colour_data = 24'b001010101100010100011000;
		13'b1001001001000: colour_data = 24'b111111110000000010010110;
		13'b1001001001001: colour_data = 24'b111111110000000010010110;
		13'b1001001001010: colour_data = 24'b111111110000000010010110;
		13'b1001001001011: colour_data = 24'b111111110000000010010110;
		13'b1001001001100: colour_data = 24'b000110000101000100011000;
		13'b1001001001101: colour_data = 24'b111111110000000010010110;
		13'b1001001001110: colour_data = 24'b111111110000000010010110;
		13'b1001001001111: colour_data = 24'b111111110000000010010110;
		13'b1001001010000: colour_data = 24'b000110000110110100011000;
		13'b1001001010001: colour_data = 24'b111111110000000010010110;
		13'b1001001010010: colour_data = 24'b111111110000000010010110;
		13'b1001001010011: colour_data = 24'b111111110000000010010110;
		13'b1001001010100: colour_data = 24'b111111110000000010010110;
		13'b1001001010101: colour_data = 24'b000110000110110100011000;
		13'b1001001010110: colour_data = 24'b111111110000000010010110;
		13'b1001001010111: colour_data = 24'b111111110000000010010110;
		13'b1001001011000: colour_data = 24'b111111110000000010010110;
		13'b1001001011001: colour_data = 24'b111111110000000010010110;
		13'b1001001011010: colour_data = 24'b001010101100010100011000;
		13'b1001001011011: colour_data = 24'b111111110000000010010110;
		13'b1001001011100: colour_data = 24'b111111110000000010010110;
		13'b1001001011101: colour_data = 24'b111111110000000010010110;
		13'b1001001011110: colour_data = 24'b000110000110110100011000;
		13'b1001001011111: colour_data = 24'b000110000101000100011000;
		13'b1001001100000: colour_data = 24'b111111110000000010010110;
		13'b1001001100001: colour_data = 24'b111111110000000010010110;
		13'b1001001100010: colour_data = 24'b111111110000000010010110;
		13'b1001001100011: colour_data = 24'b000110000110110100011000;
		13'b1001001100100: colour_data = 24'b111111110000000010010110;
		13'b1001001100101: colour_data = 24'b111111110000000010010110;
		13'b1001001100110: colour_data = 24'b111111110000000010010110;
		13'b1001001100111: colour_data = 24'b111111110000000010010110;
		13'b1001001101000: colour_data = 24'b000110000110110100011000;
		13'b1001001101001: colour_data = 24'b111111110000000010010110;
		13'b1001001101010: colour_data = 24'b111111110000000010010110;
		13'b1001001101011: colour_data = 24'b111111110000000010010110;
		13'b1001001101100: colour_data = 24'b111111110000000010010110;
		13'b1001001101101: colour_data = 24'b001010101100010100011000;
		13'b1001001101110: colour_data = 24'b111111110000000010010110;
		13'b1001001101111: colour_data = 24'b111111110000000010010110;
		13'b1001001110000: colour_data = 24'b111111110000000010010110;
		13'b1001001110001: colour_data = 24'b000110000110110100011000;
		13'b1001001110010: colour_data = 24'b000110000101000100011000;
		13'b1001001110011: colour_data = 24'b111111110000000010010110;
		13'b1001001110100: colour_data = 24'b111111110000000010010110;
		13'b1001001110101: colour_data = 24'b111111110000000010010110;
		13'b1001001110110: colour_data = 24'b000110000110110100011000;
		13'b1001001110111: colour_data = 24'b111111110000000010010110;
		13'b1001001111000: colour_data = 24'b111111110000000010010110;
		13'b1001001111001: colour_data = 24'b111111110000000010010110;
		13'b1001001111010: colour_data = 24'b111111110000000010010110;
		13'b1001001111011: colour_data = 24'b001010101100010100011000;
		13'b1001001111100: colour_data = 24'b111111110000000010010110;
		13'b1001001111101: colour_data = 24'b111111110000000010010110;
		13'b1001001111110: colour_data = 24'b111111110000000010010110;
		13'b1001001111111: colour_data = 24'b111111110000000010010110;
		13'b1001010000000: colour_data = 24'b000110000101000100011000;
		13'b1001010000001: colour_data = 24'b111111110000000010010110;
		13'b1001010000010: colour_data = 24'b111111110000000010010110;
		13'b1001010000011: colour_data = 24'b111111110000000010010110;
		13'b1001010000100: colour_data = 24'b000110000110110100011000;
		13'b1001010000101: colour_data = 24'b001010101100010100011000;
		13'b1001010000110: colour_data = 24'b111111110000000010010110;
		13'b1001010000111: colour_data = 24'b111111110000000010010110;
		13'b1001010001000: colour_data = 24'b111111110000000010010110;
		13'b1001010001001: colour_data = 24'b111111110000000010010110;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule