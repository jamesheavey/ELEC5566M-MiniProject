module numbers_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [2:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [2:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		10'b0000000000: colour_data = 24'b000000000000000000000000;
		10'b0000000001: colour_data = 24'b000000000000000000000000;
		10'b0000000010: colour_data = 24'b000000000000000000000000;
		10'b0000000011: colour_data = 24'b000000000000000000000000;
		10'b0000000100: colour_data = 24'b000000000000000000000000;
		10'b0000000101: colour_data = 24'b000000000000000000000000;
		10'b0000000110: colour_data = 24'b000000000000000000000000;

		10'b0000001000: colour_data = 24'b000000000000000000000000;
		10'b0000001001: colour_data = 24'b111111111111111111111111;
		10'b0000001010: colour_data = 24'b111111111111111111111111;
		10'b0000001011: colour_data = 24'b111111111111111111111111;
		10'b0000001100: colour_data = 24'b111111111111111111111111;
		10'b0000001101: colour_data = 24'b111111111111111111111111;
		10'b0000001110: colour_data = 24'b000000000000000000000000;

		10'b0000010000: colour_data = 24'b000000000000000000000000;
		10'b0000010001: colour_data = 24'b111111111111111111111111;
		10'b0000010010: colour_data = 24'b111111111111111111111111;
		10'b0000010011: colour_data = 24'b111111111111111111111111;
		10'b0000010100: colour_data = 24'b111111111111111111111111;
		10'b0000010101: colour_data = 24'b111111111111111111111111;
		10'b0000010110: colour_data = 24'b000000000000000000000000;

		10'b0000011000: colour_data = 24'b000000000000000000000000;
		10'b0000011001: colour_data = 24'b111111111111111111111111;
		10'b0000011010: colour_data = 24'b111111111111111111111111;
		10'b0000011011: colour_data = 24'b000000000000000000000000;
		10'b0000011100: colour_data = 24'b111111111111111111111111;
		10'b0000011101: colour_data = 24'b111111111111111111111111;
		10'b0000011110: colour_data = 24'b000000000000000000000000;

		10'b0000100000: colour_data = 24'b000000000000000000000000;
		10'b0000100001: colour_data = 24'b111111111111111111111111;
		10'b0000100010: colour_data = 24'b111111111111111111111111;
		10'b0000100011: colour_data = 24'b000000000000000000000000;
		10'b0000100100: colour_data = 24'b111111111111111111111111;
		10'b0000100101: colour_data = 24'b111111111111111111111111;
		10'b0000100110: colour_data = 24'b000000000000000000000000;

		10'b0000101000: colour_data = 24'b000000000000000000000000;
		10'b0000101001: colour_data = 24'b111111111111111111111111;
		10'b0000101010: colour_data = 24'b111111111111111111111111;
		10'b0000101011: colour_data = 24'b000000000000000000000000;
		10'b0000101100: colour_data = 24'b111111111111111111111111;
		10'b0000101101: colour_data = 24'b111111111111111111111111;
		10'b0000101110: colour_data = 24'b000000000000000000000000;

		10'b0000110000: colour_data = 24'b000000000000000000000000;
		10'b0000110001: colour_data = 24'b111111111111111111111111;
		10'b0000110010: colour_data = 24'b111111111111111111111111;
		10'b0000110011: colour_data = 24'b000000000000000000000000;
		10'b0000110100: colour_data = 24'b111111111111111111111111;
		10'b0000110101: colour_data = 24'b111111111111111111111111;
		10'b0000110110: colour_data = 24'b000000000000000000000000;

		10'b0000111000: colour_data = 24'b000000000000000000000000;
		10'b0000111001: colour_data = 24'b111111111111111111111111;
		10'b0000111010: colour_data = 24'b111111111111111111111111;
		10'b0000111011: colour_data = 24'b111111111111111111111111;
		10'b0000111100: colour_data = 24'b111111111111111111111111;
		10'b0000111101: colour_data = 24'b111111111111111111111111;
		10'b0000111110: colour_data = 24'b000000000000000000000000;

		10'b0001000000: colour_data = 24'b000000000000000000000000;
		10'b0001000001: colour_data = 24'b111111111111111111111111;
		10'b0001000010: colour_data = 24'b111111111111111111111111;
		10'b0001000011: colour_data = 24'b111111111111111111111111;
		10'b0001000100: colour_data = 24'b111111111111111111111111;
		10'b0001000101: colour_data = 24'b111111111111111111111111;
		10'b0001000110: colour_data = 24'b000000000000000000000000;

		10'b0001001000: colour_data = 24'b000000000000000000000000;
		10'b0001001001: colour_data = 24'b000000000000000000000000;
		10'b0001001010: colour_data = 24'b000000000000000000000000;
		10'b0001001011: colour_data = 24'b000000000000000000000000;
		10'b0001001100: colour_data = 24'b000000000000000000000000;
		10'b0001001101: colour_data = 24'b000000000000000000000000;
		10'b0001001110: colour_data = 24'b000000000000000000000000;

		10'b0001010000: colour_data = 24'b111111110000000010010110;
		10'b0001010001: colour_data = 24'b000000000000000000000000;
		10'b0001010010: colour_data = 24'b000000000000000000000000;
		10'b0001010011: colour_data = 24'b000000000000000000000000;
		10'b0001010100: colour_data = 24'b000000000000000000000000;
		10'b0001010101: colour_data = 24'b000000000000000000000000;
		10'b0001010110: colour_data = 24'b111111110000000010010110;

		10'b0001011000: colour_data = 24'b111111110000000010010110;
		10'b0001011001: colour_data = 24'b000000000000000000000000;
		10'b0001011010: colour_data = 24'b111111111111111111111111;
		10'b0001011011: colour_data = 24'b111111111111111111111111;
		10'b0001011100: colour_data = 24'b111111111111111111111111;
		10'b0001011101: colour_data = 24'b000000000000000000000000;
		10'b0001011110: colour_data = 24'b111111110000000010010110;

		10'b0001100000: colour_data = 24'b111111110000000010010110;
		10'b0001100001: colour_data = 24'b000000000000000000000000;
		10'b0001100010: colour_data = 24'b111111111111111111111111;
		10'b0001100011: colour_data = 24'b111111111111111111111111;
		10'b0001100100: colour_data = 24'b111111111111111111111111;
		10'b0001100101: colour_data = 24'b000000000000000000000000;
		10'b0001100110: colour_data = 24'b111111110000000010010110;

		10'b0001101000: colour_data = 24'b111111110000000010010110;
		10'b0001101001: colour_data = 24'b000000000000000000000000;
		10'b0001101010: colour_data = 24'b000000000000000000000000;
		10'b0001101011: colour_data = 24'b111111111111111111111111;
		10'b0001101100: colour_data = 24'b111111111111111111111111;
		10'b0001101101: colour_data = 24'b000000000000000000000000;
		10'b0001101110: colour_data = 24'b111111110000000010010110;

		10'b0001110000: colour_data = 24'b111111110000000010010110;
		10'b0001110001: colour_data = 24'b111111110000000010010110;
		10'b0001110010: colour_data = 24'b000000000000000000000000;
		10'b0001110011: colour_data = 24'b111111111111111111111111;
		10'b0001110100: colour_data = 24'b111111111111111111111111;
		10'b0001110101: colour_data = 24'b000000000000000000000000;
		10'b0001110110: colour_data = 24'b111111110000000010010110;

		10'b0001111000: colour_data = 24'b111111110000000010010110;
		10'b0001111001: colour_data = 24'b111111110000000010010110;
		10'b0001111010: colour_data = 24'b000000000000000000000000;
		10'b0001111011: colour_data = 24'b111111111111111111111111;
		10'b0001111100: colour_data = 24'b111111111111111111111111;
		10'b0001111101: colour_data = 24'b000000000000000000000000;
		10'b0001111110: colour_data = 24'b111111110000000010010110;

		10'b0010000000: colour_data = 24'b111111110000000010010110;
		10'b0010000001: colour_data = 24'b111111110000000010010110;
		10'b0010000010: colour_data = 24'b000000000000000000000000;
		10'b0010000011: colour_data = 24'b111111111111111111111111;
		10'b0010000100: colour_data = 24'b111111111111111111111111;
		10'b0010000101: colour_data = 24'b000000000000000000000000;
		10'b0010000110: colour_data = 24'b111111110000000010010110;

		10'b0010001000: colour_data = 24'b111111110000000010010110;
		10'b0010001001: colour_data = 24'b111111110000000010010110;
		10'b0010001010: colour_data = 24'b000000000000000000000000;
		10'b0010001011: colour_data = 24'b111111111111111111111111;
		10'b0010001100: colour_data = 24'b111111111111111111111111;
		10'b0010001101: colour_data = 24'b000000000000000000000000;
		10'b0010001110: colour_data = 24'b111111110000000010010110;

		10'b0010010000: colour_data = 24'b111111110000000010010110;
		10'b0010010001: colour_data = 24'b111111110000000010010110;
		10'b0010010010: colour_data = 24'b000000000000000000000000;
		10'b0010010011: colour_data = 24'b111111111111111111111111;
		10'b0010010100: colour_data = 24'b111111111111111111111111;
		10'b0010010101: colour_data = 24'b000000000000000000000000;
		10'b0010010110: colour_data = 24'b111111110000000010010110;

		10'b0010011000: colour_data = 24'b111111110000000010010110;
		10'b0010011001: colour_data = 24'b111111110000000010010110;
		10'b0010011010: colour_data = 24'b000000000000000000000000;
		10'b0010011011: colour_data = 24'b000000000000000000000000;
		10'b0010011100: colour_data = 24'b000000000000000000000000;
		10'b0010011101: colour_data = 24'b000000000000000000000000;
		10'b0010011110: colour_data = 24'b111111110000000010010110;

		10'b0010100000: colour_data = 24'b000000000000000000000000;
		10'b0010100001: colour_data = 24'b000000000000000000000000;
		10'b0010100010: colour_data = 24'b000000000000000000000000;
		10'b0010100011: colour_data = 24'b000000000000000000000000;
		10'b0010100100: colour_data = 24'b000000000000000000000000;
		10'b0010100101: colour_data = 24'b000000000000000000000000;
		10'b0010100110: colour_data = 24'b000000000000000000000000;

		10'b0010101000: colour_data = 24'b000000000000000000000000;
		10'b0010101001: colour_data = 24'b111111111111111111111111;
		10'b0010101010: colour_data = 24'b111111111111111111111111;
		10'b0010101011: colour_data = 24'b111111111111111111111111;
		10'b0010101100: colour_data = 24'b111111111111111111111111;
		10'b0010101101: colour_data = 24'b111111111111111111111111;
		10'b0010101110: colour_data = 24'b000000000000000000000000;

		10'b0010110000: colour_data = 24'b000000000000000000000000;
		10'b0010110001: colour_data = 24'b111111111111111111111111;
		10'b0010110010: colour_data = 24'b111111111111111111111111;
		10'b0010110011: colour_data = 24'b111111111111111111111111;
		10'b0010110100: colour_data = 24'b111111111111111111111111;
		10'b0010110101: colour_data = 24'b111111111111111111111111;
		10'b0010110110: colour_data = 24'b000000000000000000000000;

		10'b0010111000: colour_data = 24'b000000000000000000000000;
		10'b0010111001: colour_data = 24'b000000000000000000000000;
		10'b0010111010: colour_data = 24'b000000000000000000000000;
		10'b0010111011: colour_data = 24'b000000000000000000000000;
		10'b0010111100: colour_data = 24'b111111111111111111111111;
		10'b0010111101: colour_data = 24'b111111111111111111111111;
		10'b0010111110: colour_data = 24'b000000000000000000000000;

		10'b0011000000: colour_data = 24'b000000000000000000000000;
		10'b0011000001: colour_data = 24'b111111111111111111111111;
		10'b0011000010: colour_data = 24'b111111111111111111111111;
		10'b0011000011: colour_data = 24'b111111111111111111111111;
		10'b0011000100: colour_data = 24'b111111111111111111111111;
		10'b0011000101: colour_data = 24'b111111111111111111111111;
		10'b0011000110: colour_data = 24'b000000000000000000000000;

		10'b0011001000: colour_data = 24'b000000000000000000000000;
		10'b0011001001: colour_data = 24'b111111111111111111111111;
		10'b0011001010: colour_data = 24'b111111111111111111111111;
		10'b0011001011: colour_data = 24'b111111111111111111111111;
		10'b0011001100: colour_data = 24'b111111111111111111111111;
		10'b0011001101: colour_data = 24'b111111111111111111111111;
		10'b0011001110: colour_data = 24'b000000000000000000000000;

		10'b0011010000: colour_data = 24'b000000000000000000000000;
		10'b0011010001: colour_data = 24'b111111111111111111111111;
		10'b0011010010: colour_data = 24'b111111111111111111111111;
		10'b0011010011: colour_data = 24'b000000000000000000000000;
		10'b0011010100: colour_data = 24'b000000000000000000000000;
		10'b0011010101: colour_data = 24'b000000000000000000000000;
		10'b0011010110: colour_data = 24'b000000000000000000000000;

		10'b0011011000: colour_data = 24'b000000000000000000000000;
		10'b0011011001: colour_data = 24'b111111111111111111111111;
		10'b0011011010: colour_data = 24'b111111111111111111111111;
		10'b0011011011: colour_data = 24'b111111111111111111111111;
		10'b0011011100: colour_data = 24'b111111111111111111111111;
		10'b0011011101: colour_data = 24'b111111111111111111111111;
		10'b0011011110: colour_data = 24'b000000000000000000000000;

		10'b0011100000: colour_data = 24'b000000000000000000000000;
		10'b0011100001: colour_data = 24'b111111111111111111111111;
		10'b0011100010: colour_data = 24'b111111111111111111111111;
		10'b0011100011: colour_data = 24'b111111111111111111111111;
		10'b0011100100: colour_data = 24'b111111111111111111111111;
		10'b0011100101: colour_data = 24'b111111111111111111111111;
		10'b0011100110: colour_data = 24'b000000000000000000000000;

		10'b0011101000: colour_data = 24'b000000000000000000000000;
		10'b0011101001: colour_data = 24'b000000000000000000000000;
		10'b0011101010: colour_data = 24'b000000000000000000000000;
		10'b0011101011: colour_data = 24'b000000000000000000000000;
		10'b0011101100: colour_data = 24'b000000000000000000000000;
		10'b0011101101: colour_data = 24'b000000000000000000000000;
		10'b0011101110: colour_data = 24'b000000000000000000000000;

		10'b0011110000: colour_data = 24'b000000000000000000000000;
		10'b0011110001: colour_data = 24'b000000000000000000000000;
		10'b0011110010: colour_data = 24'b000000000000000000000000;
		10'b0011110011: colour_data = 24'b000000000000000000000000;
		10'b0011110100: colour_data = 24'b000000000000000000000000;
		10'b0011110101: colour_data = 24'b000000000000000000000000;
		10'b0011110110: colour_data = 24'b000000000000000000000000;

		10'b0011111000: colour_data = 24'b000000000000000000000000;
		10'b0011111001: colour_data = 24'b111111111111111111111111;
		10'b0011111010: colour_data = 24'b111111111111111111111111;
		10'b0011111011: colour_data = 24'b111111111111111111111111;
		10'b0011111100: colour_data = 24'b111111111111111111111111;
		10'b0011111101: colour_data = 24'b111111111111111111111111;
		10'b0011111110: colour_data = 24'b000000000000000000000000;

		10'b0100000000: colour_data = 24'b000000000000000000000000;
		10'b0100000001: colour_data = 24'b111111111111111111111111;
		10'b0100000010: colour_data = 24'b111111111111111111111111;
		10'b0100000011: colour_data = 24'b111111111111111111111111;
		10'b0100000100: colour_data = 24'b111111111111111111111111;
		10'b0100000101: colour_data = 24'b111111111111111111111111;
		10'b0100000110: colour_data = 24'b000000000000000000000000;

		10'b0100001000: colour_data = 24'b000000000000000000000000;
		10'b0100001001: colour_data = 24'b000000000000000000000000;
		10'b0100001010: colour_data = 24'b000000000000000000000000;
		10'b0100001011: colour_data = 24'b000000000000000000000000;
		10'b0100001100: colour_data = 24'b111111111111111111111111;
		10'b0100001101: colour_data = 24'b111111111111111111111111;
		10'b0100001110: colour_data = 24'b000000000000000000000000;

		10'b0100010000: colour_data = 24'b000000000000000000000000;
		10'b0100010001: colour_data = 24'b111111111111111111111111;
		10'b0100010010: colour_data = 24'b111111111111111111111111;
		10'b0100010011: colour_data = 24'b111111111111111111111111;
		10'b0100010100: colour_data = 24'b111111111111111111111111;
		10'b0100010101: colour_data = 24'b111111111111111111111111;
		10'b0100010110: colour_data = 24'b000000000000000000000000;

		10'b0100011000: colour_data = 24'b000000000000000000000000;
		10'b0100011001: colour_data = 24'b111111111111111111111111;
		10'b0100011010: colour_data = 24'b111111111111111111111111;
		10'b0100011011: colour_data = 24'b111111111111111111111111;
		10'b0100011100: colour_data = 24'b111111111111111111111111;
		10'b0100011101: colour_data = 24'b111111111111111111111111;
		10'b0100011110: colour_data = 24'b000000000000000000000000;

		10'b0100100000: colour_data = 24'b000000000000000000000000;
		10'b0100100001: colour_data = 24'b000000000000000000000000;
		10'b0100100010: colour_data = 24'b000000000000000000000000;
		10'b0100100011: colour_data = 24'b000000000000000000000000;
		10'b0100100100: colour_data = 24'b111111111111111111111111;
		10'b0100100101: colour_data = 24'b111111111111111111111111;
		10'b0100100110: colour_data = 24'b000000000000000000000000;

		10'b0100101000: colour_data = 24'b000000000000000000000000;
		10'b0100101001: colour_data = 24'b111111111111111111111111;
		10'b0100101010: colour_data = 24'b111111111111111111111111;
		10'b0100101011: colour_data = 24'b111111111111111111111111;
		10'b0100101100: colour_data = 24'b111111111111111111111111;
		10'b0100101101: colour_data = 24'b111111111111111111111111;
		10'b0100101110: colour_data = 24'b000000000000000000000000;

		10'b0100110000: colour_data = 24'b000000000000000000000000;
		10'b0100110001: colour_data = 24'b111111111111111111111111;
		10'b0100110010: colour_data = 24'b111111111111111111111111;
		10'b0100110011: colour_data = 24'b111111111111111111111111;
		10'b0100110100: colour_data = 24'b111111111111111111111111;
		10'b0100110101: colour_data = 24'b111111111111111111111111;
		10'b0100110110: colour_data = 24'b000000000000000000000000;

		10'b0100111000: colour_data = 24'b000000000000000000000000;
		10'b0100111001: colour_data = 24'b000000000000000000000000;
		10'b0100111010: colour_data = 24'b000000000000000000000000;
		10'b0100111011: colour_data = 24'b000000000000000000000000;
		10'b0100111100: colour_data = 24'b000000000000000000000000;
		10'b0100111101: colour_data = 24'b000000000000000000000000;
		10'b0100111110: colour_data = 24'b000000000000000000000000;

		10'b0101000000: colour_data = 24'b000000000000000000000000;
		10'b0101000001: colour_data = 24'b000000000000000000000000;
		10'b0101000010: colour_data = 24'b000000000000000000000000;
		10'b0101000011: colour_data = 24'b000000000000000000000000;
		10'b0101000100: colour_data = 24'b000000000000000000000000;
		10'b0101000101: colour_data = 24'b000000000000000000000000;
		10'b0101000110: colour_data = 24'b000000000000000000000000;

		10'b0101001000: colour_data = 24'b000000000000000000000000;
		10'b0101001001: colour_data = 24'b111111111111111111111111;
		10'b0101001010: colour_data = 24'b111111111111111111111111;
		10'b0101001011: colour_data = 24'b000000000000000000000000;
		10'b0101001100: colour_data = 24'b111111111111111111111111;
		10'b0101001101: colour_data = 24'b111111111111111111111111;
		10'b0101001110: colour_data = 24'b000000000000000000000000;

		10'b0101010000: colour_data = 24'b000000000000000000000000;
		10'b0101010001: colour_data = 24'b111111111111111111111111;
		10'b0101010010: colour_data = 24'b111111111111111111111111;
		10'b0101010011: colour_data = 24'b000000000000000000000000;
		10'b0101010100: colour_data = 24'b111111111111111111111111;
		10'b0101010101: colour_data = 24'b111111111111111111111111;
		10'b0101010110: colour_data = 24'b000000000000000000000000;

		10'b0101011000: colour_data = 24'b000000000000000000000000;
		10'b0101011001: colour_data = 24'b111111111111111111111111;
		10'b0101011010: colour_data = 24'b111111111111111111111111;
		10'b0101011011: colour_data = 24'b000000000000000000000000;
		10'b0101011100: colour_data = 24'b111111111111111111111111;
		10'b0101011101: colour_data = 24'b111111111111111111111111;
		10'b0101011110: colour_data = 24'b000000000000000000000000;

		10'b0101100000: colour_data = 24'b000000000000000000000000;
		10'b0101100001: colour_data = 24'b111111111111111111111111;
		10'b0101100010: colour_data = 24'b111111111111111111111111;
		10'b0101100011: colour_data = 24'b111111111111111111111111;
		10'b0101100100: colour_data = 24'b111111111111111111111111;
		10'b0101100101: colour_data = 24'b111111111111111111111111;
		10'b0101100110: colour_data = 24'b000000000000000000000000;

		10'b0101101000: colour_data = 24'b000000000000000000000000;
		10'b0101101001: colour_data = 24'b111111111111111111111111;
		10'b0101101010: colour_data = 24'b111111111111111111111111;
		10'b0101101011: colour_data = 24'b111111111111111111111111;
		10'b0101101100: colour_data = 24'b111111111111111111111111;
		10'b0101101101: colour_data = 24'b111111111111111111111111;
		10'b0101101110: colour_data = 24'b000000000000000000000000;

		10'b0101110000: colour_data = 24'b000000000000000000000000;
		10'b0101110001: colour_data = 24'b000000000000000000000000;
		10'b0101110010: colour_data = 24'b000000000000000000000000;
		10'b0101110011: colour_data = 24'b000000000000000000000000;
		10'b0101110100: colour_data = 24'b111111111111111111111111;
		10'b0101110101: colour_data = 24'b111111111111111111111111;
		10'b0101110110: colour_data = 24'b000000000000000000000000;

		10'b0101111000: colour_data = 24'b111111110000000010010110;
		10'b0101111001: colour_data = 24'b111111110000000010010110;
		10'b0101111010: colour_data = 24'b111111110000000010010110;
		10'b0101111011: colour_data = 24'b000000000000000000000000;
		10'b0101111100: colour_data = 24'b111111111111111111111111;
		10'b0101111101: colour_data = 24'b111111111111111111111111;
		10'b0101111110: colour_data = 24'b000000000000000000000000;

		10'b0110000000: colour_data = 24'b111111110000000010010110;
		10'b0110000001: colour_data = 24'b111111110000000010010110;
		10'b0110000010: colour_data = 24'b111111110000000010010110;
		10'b0110000011: colour_data = 24'b000000000000000000000000;
		10'b0110000100: colour_data = 24'b111111111111111111111111;
		10'b0110000101: colour_data = 24'b111111111111111111111111;
		10'b0110000110: colour_data = 24'b000000000000000000000000;

		10'b0110001000: colour_data = 24'b111111110000000010010110;
		10'b0110001001: colour_data = 24'b111111110000000010010110;
		10'b0110001010: colour_data = 24'b111111110000000010010110;
		10'b0110001011: colour_data = 24'b000000000000000000000000;
		10'b0110001100: colour_data = 24'b000000000000000000000000;
		10'b0110001101: colour_data = 24'b000000000000000000000000;
		10'b0110001110: colour_data = 24'b000000000000000000000000;

		10'b0110010000: colour_data = 24'b000000000000000000000000;
		10'b0110010001: colour_data = 24'b000000000000000000000000;
		10'b0110010010: colour_data = 24'b000000000000000000000000;
		10'b0110010011: colour_data = 24'b000000000000000000000000;
		10'b0110010100: colour_data = 24'b000000000000000000000000;
		10'b0110010101: colour_data = 24'b000000000000000000000000;
		10'b0110010110: colour_data = 24'b000000000000000000000000;

		10'b0110011000: colour_data = 24'b000000000000000000000000;
		10'b0110011001: colour_data = 24'b111111111111111111111111;
		10'b0110011010: colour_data = 24'b111111111111111111111111;
		10'b0110011011: colour_data = 24'b111111111111111111111111;
		10'b0110011100: colour_data = 24'b111111111111111111111111;
		10'b0110011101: colour_data = 24'b111111111111111111111111;
		10'b0110011110: colour_data = 24'b000000000000000000000000;

		10'b0110100000: colour_data = 24'b000000000000000000000000;
		10'b0110100001: colour_data = 24'b111111111111111111111111;
		10'b0110100010: colour_data = 24'b111111111111111111111111;
		10'b0110100011: colour_data = 24'b111111111111111111111111;
		10'b0110100100: colour_data = 24'b111111111111111111111111;
		10'b0110100101: colour_data = 24'b111111111111111111111111;
		10'b0110100110: colour_data = 24'b000000000000000000000000;

		10'b0110101000: colour_data = 24'b000000000000000000000000;
		10'b0110101001: colour_data = 24'b111111111111111111111111;
		10'b0110101010: colour_data = 24'b111111111111111111111111;
		10'b0110101011: colour_data = 24'b000000000000000000000000;
		10'b0110101100: colour_data = 24'b000000000000000000000000;
		10'b0110101101: colour_data = 24'b000000000000000000000000;
		10'b0110101110: colour_data = 24'b000000000000000000000000;

		10'b0110110000: colour_data = 24'b000000000000000000000000;
		10'b0110110001: colour_data = 24'b111111111111111111111111;
		10'b0110110010: colour_data = 24'b111111111111111111111111;
		10'b0110110011: colour_data = 24'b111111111111111111111111;
		10'b0110110100: colour_data = 24'b111111111111111111111111;
		10'b0110110101: colour_data = 24'b111111111111111111111111;
		10'b0110110110: colour_data = 24'b000000000000000000000000;

		10'b0110111000: colour_data = 24'b000000000000000000000000;
		10'b0110111001: colour_data = 24'b111111111111111111111111;
		10'b0110111010: colour_data = 24'b111111111111111111111111;
		10'b0110111011: colour_data = 24'b111111111111111111111111;
		10'b0110111100: colour_data = 24'b111111111111111111111111;
		10'b0110111101: colour_data = 24'b111111111111111111111111;
		10'b0110111110: colour_data = 24'b000000000000000000000000;

		10'b0111000000: colour_data = 24'b000000000000000000000000;
		10'b0111000001: colour_data = 24'b000000000000000000000000;
		10'b0111000010: colour_data = 24'b000000000000000000000000;
		10'b0111000011: colour_data = 24'b000000000000000000000000;
		10'b0111000100: colour_data = 24'b111111111111111111111111;
		10'b0111000101: colour_data = 24'b111111111111111111111111;
		10'b0111000110: colour_data = 24'b000000000000000000000000;

		10'b0111001000: colour_data = 24'b000000000000000000000000;
		10'b0111001001: colour_data = 24'b111111111111111111111111;
		10'b0111001010: colour_data = 24'b111111111111111111111111;
		10'b0111001011: colour_data = 24'b111111111111111111111111;
		10'b0111001100: colour_data = 24'b111111111111111111111111;
		10'b0111001101: colour_data = 24'b111111111111111111111111;
		10'b0111001110: colour_data = 24'b000000000000000000000000;

		10'b0111010000: colour_data = 24'b000000000000000000000000;
		10'b0111010001: colour_data = 24'b111111111111111111111111;
		10'b0111010010: colour_data = 24'b111111111111111111111111;
		10'b0111010011: colour_data = 24'b111111111111111111111111;
		10'b0111010100: colour_data = 24'b111111111111111111111111;
		10'b0111010101: colour_data = 24'b111111111111111111111111;
		10'b0111010110: colour_data = 24'b000000000000000000000000;

		10'b0111011000: colour_data = 24'b000000000000000000000000;
		10'b0111011001: colour_data = 24'b000000000000000000000000;
		10'b0111011010: colour_data = 24'b000000000000000000000000;
		10'b0111011011: colour_data = 24'b000000000000000000000000;
		10'b0111011100: colour_data = 24'b000000000000000000000000;
		10'b0111011101: colour_data = 24'b000000000000000000000000;
		10'b0111011110: colour_data = 24'b000000000000000000000000;

		10'b0111100000: colour_data = 24'b000000000000000000000000;
		10'b0111100001: colour_data = 24'b000000000000000000000000;
		10'b0111100010: colour_data = 24'b000000000000000000000000;
		10'b0111100011: colour_data = 24'b000000000000000000000000;
		10'b0111100100: colour_data = 24'b000000000000000000000000;
		10'b0111100101: colour_data = 24'b000000000000000000000000;
		10'b0111100110: colour_data = 24'b000000000000000000000000;

		10'b0111101000: colour_data = 24'b000000000000000000000000;
		10'b0111101001: colour_data = 24'b111111111111111111111111;
		10'b0111101010: colour_data = 24'b111111111111111111111111;
		10'b0111101011: colour_data = 24'b111111111111111111111111;
		10'b0111101100: colour_data = 24'b111111111111111111111111;
		10'b0111101101: colour_data = 24'b111111111111111111111111;
		10'b0111101110: colour_data = 24'b000000000000000000000000;

		10'b0111110000: colour_data = 24'b000000000000000000000000;
		10'b0111110001: colour_data = 24'b111111111111111111111111;
		10'b0111110010: colour_data = 24'b111111111111111111111111;
		10'b0111110011: colour_data = 24'b111111111111111111111111;
		10'b0111110100: colour_data = 24'b111111111111111111111111;
		10'b0111110101: colour_data = 24'b111111111111111111111111;
		10'b0111110110: colour_data = 24'b000000000000000000000000;

		10'b0111111000: colour_data = 24'b000000000000000000000000;
		10'b0111111001: colour_data = 24'b111111111111111111111111;
		10'b0111111010: colour_data = 24'b111111111111111111111111;
		10'b0111111011: colour_data = 24'b000000000000000000000000;
		10'b0111111100: colour_data = 24'b000000000000000000000000;
		10'b0111111101: colour_data = 24'b000000000000000000000000;
		10'b0111111110: colour_data = 24'b000000000000000000000000;

		10'b1000000000: colour_data = 24'b000000000000000000000000;
		10'b1000000001: colour_data = 24'b111111111111111111111111;
		10'b1000000010: colour_data = 24'b111111111111111111111111;
		10'b1000000011: colour_data = 24'b111111111111111111111111;
		10'b1000000100: colour_data = 24'b111111111111111111111111;
		10'b1000000101: colour_data = 24'b111111111111111111111111;
		10'b1000000110: colour_data = 24'b000000000000000000000000;

		10'b1000001000: colour_data = 24'b000000000000000000000000;
		10'b1000001001: colour_data = 24'b111111111111111111111111;
		10'b1000001010: colour_data = 24'b111111111111111111111111;
		10'b1000001011: colour_data = 24'b111111111111111111111111;
		10'b1000001100: colour_data = 24'b111111111111111111111111;
		10'b1000001101: colour_data = 24'b111111111111111111111111;
		10'b1000001110: colour_data = 24'b000000000000000000000000;

		10'b1000010000: colour_data = 24'b000000000000000000000000;
		10'b1000010001: colour_data = 24'b111111111111111111111111;
		10'b1000010010: colour_data = 24'b111111111111111111111111;
		10'b1000010011: colour_data = 24'b000000000000000000000000;
		10'b1000010100: colour_data = 24'b111111111111111111111111;
		10'b1000010101: colour_data = 24'b111111111111111111111111;
		10'b1000010110: colour_data = 24'b000000000000000000000000;

		10'b1000011000: colour_data = 24'b000000000000000000000000;
		10'b1000011001: colour_data = 24'b111111111111111111111111;
		10'b1000011010: colour_data = 24'b111111111111111111111111;
		10'b1000011011: colour_data = 24'b111111111111111111111111;
		10'b1000011100: colour_data = 24'b111111111111111111111111;
		10'b1000011101: colour_data = 24'b111111111111111111111111;
		10'b1000011110: colour_data = 24'b000000000000000000000000;

		10'b1000100000: colour_data = 24'b000000000000000000000000;
		10'b1000100001: colour_data = 24'b111111111111111111111111;
		10'b1000100010: colour_data = 24'b111111111111111111111111;
		10'b1000100011: colour_data = 24'b111111111111111111111111;
		10'b1000100100: colour_data = 24'b111111111111111111111111;
		10'b1000100101: colour_data = 24'b111111111111111111111111;
		10'b1000100110: colour_data = 24'b000000000000000000000000;

		10'b1000101000: colour_data = 24'b000000000000000000000000;
		10'b1000101001: colour_data = 24'b000000000000000000000000;
		10'b1000101010: colour_data = 24'b000000000000000000000000;
		10'b1000101011: colour_data = 24'b000000000000000000000000;
		10'b1000101100: colour_data = 24'b000000000000000000000000;
		10'b1000101101: colour_data = 24'b000000000000000000000000;
		10'b1000101110: colour_data = 24'b000000000000000000000000;

		10'b1000110000: colour_data = 24'b000000000000000000000000;
		10'b1000110001: colour_data = 24'b000000000000000000000000;
		10'b1000110010: colour_data = 24'b000000000000000000000000;
		10'b1000110011: colour_data = 24'b000000000000000000000000;
		10'b1000110100: colour_data = 24'b000000000000000000000000;
		10'b1000110101: colour_data = 24'b000000000000000000000000;
		10'b1000110110: colour_data = 24'b000000000000000000000000;

		10'b1000111000: colour_data = 24'b000000000000000000000000;
		10'b1000111001: colour_data = 24'b111111111111111111111111;
		10'b1000111010: colour_data = 24'b111111111111111111111111;
		10'b1000111011: colour_data = 24'b111111111111111111111111;
		10'b1000111100: colour_data = 24'b111111111111111111111111;
		10'b1000111101: colour_data = 24'b111111111111111111111111;
		10'b1000111110: colour_data = 24'b000000000000000000000000;

		10'b1001000000: colour_data = 24'b000000000000000000000000;
		10'b1001000001: colour_data = 24'b111111111111111111111111;
		10'b1001000010: colour_data = 24'b111111111111111111111111;
		10'b1001000011: colour_data = 24'b111111111111111111111111;
		10'b1001000100: colour_data = 24'b111111111111111111111111;
		10'b1001000101: colour_data = 24'b111111111111111111111111;
		10'b1001000110: colour_data = 24'b000000000000000000000000;

		10'b1001001000: colour_data = 24'b000000000000000000000000;
		10'b1001001001: colour_data = 24'b000000000000000000000000;
		10'b1001001010: colour_data = 24'b000000000000000000000000;
		10'b1001001011: colour_data = 24'b000000000000000000000000;
		10'b1001001100: colour_data = 24'b111111111111111111111111;
		10'b1001001101: colour_data = 24'b111111111111111111111111;
		10'b1001001110: colour_data = 24'b000000000000000000000000;

		10'b1001010000: colour_data = 24'b111111110000000010010110;
		10'b1001010001: colour_data = 24'b111111110000000010010110;
		10'b1001010010: colour_data = 24'b111111110000000010010110;
		10'b1001010011: colour_data = 24'b000000000000000000000000;
		10'b1001010100: colour_data = 24'b111111111111111111111111;
		10'b1001010101: colour_data = 24'b111111111111111111111111;
		10'b1001010110: colour_data = 24'b000000000000000000000000;

		10'b1001011000: colour_data = 24'b111111110000000010010110;
		10'b1001011001: colour_data = 24'b111111110000000010010110;
		10'b1001011010: colour_data = 24'b111111110000000010010110;
		10'b1001011011: colour_data = 24'b000000000000000000000000;
		10'b1001011100: colour_data = 24'b111111111111111111111111;
		10'b1001011101: colour_data = 24'b111111111111111111111111;
		10'b1001011110: colour_data = 24'b000000000000000000000000;

		10'b1001100000: colour_data = 24'b111111110000000010010110;
		10'b1001100001: colour_data = 24'b111111110000000010010110;
		10'b1001100010: colour_data = 24'b111111110000000010010110;
		10'b1001100011: colour_data = 24'b000000000000000000000000;
		10'b1001100100: colour_data = 24'b111111111111111111111111;
		10'b1001100101: colour_data = 24'b111111111111111111111111;
		10'b1001100110: colour_data = 24'b000000000000000000000000;

		10'b1001101000: colour_data = 24'b111111110000000010010110;
		10'b1001101001: colour_data = 24'b111111110000000010010110;
		10'b1001101010: colour_data = 24'b111111110000000010010110;
		10'b1001101011: colour_data = 24'b000000000000000000000000;
		10'b1001101100: colour_data = 24'b111111111111111111111111;
		10'b1001101101: colour_data = 24'b111111111111111111111111;
		10'b1001101110: colour_data = 24'b000000000000000000000000;

		10'b1001110000: colour_data = 24'b111111110000000010010110;
		10'b1001110001: colour_data = 24'b111111110000000010010110;
		10'b1001110010: colour_data = 24'b111111110000000010010110;
		10'b1001110011: colour_data = 24'b000000000000000000000000;
		10'b1001110100: colour_data = 24'b111111111111111111111111;
		10'b1001110101: colour_data = 24'b111111111111111111111111;
		10'b1001110110: colour_data = 24'b000000000000000000000000;

		10'b1001111000: colour_data = 24'b111111110000000010010110;
		10'b1001111001: colour_data = 24'b111111110000000010010110;
		10'b1001111010: colour_data = 24'b111111110000000010010110;
		10'b1001111011: colour_data = 24'b000000000000000000000000;
		10'b1001111100: colour_data = 24'b000000000000000000000000;
		10'b1001111101: colour_data = 24'b000000000000000000000000;
		10'b1001111110: colour_data = 24'b000000000000000000000000;

		10'b1010000000: colour_data = 24'b000000000000000000000000;
		10'b1010000001: colour_data = 24'b000000000000000000000000;
		10'b1010000010: colour_data = 24'b000000000000000000000000;
		10'b1010000011: colour_data = 24'b000000000000000000000000;
		10'b1010000100: colour_data = 24'b000000000000000000000000;
		10'b1010000101: colour_data = 24'b000000000000000000000000;
		10'b1010000110: colour_data = 24'b000000000000000000000000;

		10'b1010001000: colour_data = 24'b000000000000000000000000;
		10'b1010001001: colour_data = 24'b111111111111111111111111;
		10'b1010001010: colour_data = 24'b111111111111111111111111;
		10'b1010001011: colour_data = 24'b111111111111111111111111;
		10'b1010001100: colour_data = 24'b111111111111111111111111;
		10'b1010001101: colour_data = 24'b111111111111111111111111;
		10'b1010001110: colour_data = 24'b000000000000000000000000;

		10'b1010010000: colour_data = 24'b000000000000000000000000;
		10'b1010010001: colour_data = 24'b111111111111111111111111;
		10'b1010010010: colour_data = 24'b111111111111111111111111;
		10'b1010010011: colour_data = 24'b111111111111111111111111;
		10'b1010010100: colour_data = 24'b111111111111111111111111;
		10'b1010010101: colour_data = 24'b111111111111111111111111;
		10'b1010010110: colour_data = 24'b000000000000000000000000;

		10'b1010011000: colour_data = 24'b000000000000000000000000;
		10'b1010011001: colour_data = 24'b111111111111111111111111;
		10'b1010011010: colour_data = 24'b111111111111111111111111;
		10'b1010011011: colour_data = 24'b000000000000000000000000;
		10'b1010011100: colour_data = 24'b111111111111111111111111;
		10'b1010011101: colour_data = 24'b111111111111111111111111;
		10'b1010011110: colour_data = 24'b000000000000000000000000;

		10'b1010100000: colour_data = 24'b000000000000000000000000;
		10'b1010100001: colour_data = 24'b111111111111111111111111;
		10'b1010100010: colour_data = 24'b111111111111111111111111;
		10'b1010100011: colour_data = 24'b111111111111111111111111;
		10'b1010100100: colour_data = 24'b111111111111111111111111;
		10'b1010100101: colour_data = 24'b111111111111111111111111;
		10'b1010100110: colour_data = 24'b000000000000000000000000;

		10'b1010101000: colour_data = 24'b000000000000000000000000;
		10'b1010101001: colour_data = 24'b111111111111111111111111;
		10'b1010101010: colour_data = 24'b111111111111111111111111;
		10'b1010101011: colour_data = 24'b111111111111111111111111;
		10'b1010101100: colour_data = 24'b111111111111111111111111;
		10'b1010101101: colour_data = 24'b111111111111111111111111;
		10'b1010101110: colour_data = 24'b000000000000000000000000;

		10'b1010110000: colour_data = 24'b000000000000000000000000;
		10'b1010110001: colour_data = 24'b111111111111111111111111;
		10'b1010110010: colour_data = 24'b111111111111111111111111;
		10'b1010110011: colour_data = 24'b000000000000000000000000;
		10'b1010110100: colour_data = 24'b111111111111111111111111;
		10'b1010110101: colour_data = 24'b111111111111111111111111;
		10'b1010110110: colour_data = 24'b000000000000000000000000;

		10'b1010111000: colour_data = 24'b000000000000000000000000;
		10'b1010111001: colour_data = 24'b111111111111111111111111;
		10'b1010111010: colour_data = 24'b111111111111111111111111;
		10'b1010111011: colour_data = 24'b111111111111111111111111;
		10'b1010111100: colour_data = 24'b111111111111111111111111;
		10'b1010111101: colour_data = 24'b111111111111111111111111;
		10'b1010111110: colour_data = 24'b000000000000000000000000;

		10'b1011000000: colour_data = 24'b000000000000000000000000;
		10'b1011000001: colour_data = 24'b111111111111111111111111;
		10'b1011000010: colour_data = 24'b111111111111111111111111;
		10'b1011000011: colour_data = 24'b111111111111111111111111;
		10'b1011000100: colour_data = 24'b111111111111111111111111;
		10'b1011000101: colour_data = 24'b111111111111111111111111;
		10'b1011000110: colour_data = 24'b000000000000000000000000;

		10'b1011001000: colour_data = 24'b000000000000000000000000;
		10'b1011001001: colour_data = 24'b000000000000000000000000;
		10'b1011001010: colour_data = 24'b000000000000000000000000;
		10'b1011001011: colour_data = 24'b000000000000000000000000;
		10'b1011001100: colour_data = 24'b000000000000000000000000;
		10'b1011001101: colour_data = 24'b000000000000000000000000;
		10'b1011001110: colour_data = 24'b000000000000000000000000;

		10'b1011010000: colour_data = 24'b000000000000000000000000;
		10'b1011010001: colour_data = 24'b000000000000000000000000;
		10'b1011010010: colour_data = 24'b000000000000000000000000;
		10'b1011010011: colour_data = 24'b000000000000000000000000;
		10'b1011010100: colour_data = 24'b000000000000000000000000;
		10'b1011010101: colour_data = 24'b000000000000000000000000;
		10'b1011010110: colour_data = 24'b000000000000000000000000;

		10'b1011011000: colour_data = 24'b000000000000000000000000;
		10'b1011011001: colour_data = 24'b111111111111111111111111;
		10'b1011011010: colour_data = 24'b111111111111111111111111;
		10'b1011011011: colour_data = 24'b111111111111111111111111;
		10'b1011011100: colour_data = 24'b111111111111111111111111;
		10'b1011011101: colour_data = 24'b111111111111111111111111;
		10'b1011011110: colour_data = 24'b000000000000000000000000;

		10'b1011100000: colour_data = 24'b000000000000000000000000;
		10'b1011100001: colour_data = 24'b111111111111111111111111;
		10'b1011100010: colour_data = 24'b111111111111111111111111;
		10'b1011100011: colour_data = 24'b111111111111111111111111;
		10'b1011100100: colour_data = 24'b111111111111111111111111;
		10'b1011100101: colour_data = 24'b111111111111111111111111;
		10'b1011100110: colour_data = 24'b000000000000000000000000;

		10'b1011101000: colour_data = 24'b000000000000000000000000;
		10'b1011101001: colour_data = 24'b111111111111111111111111;
		10'b1011101010: colour_data = 24'b111111111111111111111111;
		10'b1011101011: colour_data = 24'b000000000000000000000000;
		10'b1011101100: colour_data = 24'b111111111111111111111111;
		10'b1011101101: colour_data = 24'b111111111111111111111111;
		10'b1011101110: colour_data = 24'b000000000000000000000000;

		10'b1011110000: colour_data = 24'b000000000000000000000000;
		10'b1011110001: colour_data = 24'b111111111111111111111111;
		10'b1011110010: colour_data = 24'b111111111111111111111111;
		10'b1011110011: colour_data = 24'b111111111111111111111111;
		10'b1011110100: colour_data = 24'b111111111111111111111111;
		10'b1011110101: colour_data = 24'b111111111111111111111111;
		10'b1011110110: colour_data = 24'b000000000000000000000000;

		10'b1011111000: colour_data = 24'b000000000000000000000000;
		10'b1011111001: colour_data = 24'b111111111111111111111111;
		10'b1011111010: colour_data = 24'b111111111111111111111111;
		10'b1011111011: colour_data = 24'b111111111111111111111111;
		10'b1011111100: colour_data = 24'b111111111111111111111111;
		10'b1011111101: colour_data = 24'b111111111111111111111111;
		10'b1011111110: colour_data = 24'b000000000000000000000000;

		10'b1100000000: colour_data = 24'b000000000000000000000000;
		10'b1100000001: colour_data = 24'b000000000000000000000000;
		10'b1100000010: colour_data = 24'b000000000000000000000000;
		10'b1100000011: colour_data = 24'b000000000000000000000000;
		10'b1100000100: colour_data = 24'b111111111111111111111111;
		10'b1100000101: colour_data = 24'b111111111111111111111111;
		10'b1100000110: colour_data = 24'b000000000000000000000000;

		10'b1100001000: colour_data = 24'b000000000000000000000000;
		10'b1100001001: colour_data = 24'b111111111111111111111111;
		10'b1100001010: colour_data = 24'b111111111111111111111111;
		10'b1100001011: colour_data = 24'b111111111111111111111111;
		10'b1100001100: colour_data = 24'b111111111111111111111111;
		10'b1100001101: colour_data = 24'b111111111111111111111111;
		10'b1100001110: colour_data = 24'b000000000000000000000000;

		10'b1100010000: colour_data = 24'b000000000000000000000000;
		10'b1100010001: colour_data = 24'b111111111111111111111111;
		10'b1100010010: colour_data = 24'b111111111111111111111111;
		10'b1100010011: colour_data = 24'b111111111111111111111111;
		10'b1100010100: colour_data = 24'b111111111111111111111111;
		10'b1100010101: colour_data = 24'b111111111111111111111111;
		10'b1100010110: colour_data = 24'b000000000000000000000000;

		10'b1100011000: colour_data = 24'b000000000000000000000000;
		10'b1100011001: colour_data = 24'b000000000000000000000000;
		10'b1100011010: colour_data = 24'b000000000000000000000000;
		10'b1100011011: colour_data = 24'b000000000000000000000000;
		10'b1100011100: colour_data = 24'b000000000000000000000000;
		10'b1100011101: colour_data = 24'b000000000000000000000000;
		10'b1100011110: colour_data = 24'b000000000000000000000000;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule