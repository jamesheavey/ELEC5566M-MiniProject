
module bird_physics#(
	parameter BIRD_SIZE_X,
	parameter BIRD_SIZE_Y
)(
	input clk, rst, flap, 
	input [3:0] game_state,
	output reg [31:0] birdY,
	output reg [1:0] bird_state
);

localparam	START_SCREEN 	= 4'b0001,
				IN_GAME			= 4'b0010,
				PAUSE 			= 4'b0100,
				END_SCREEN 		= 4'b1000;

localparam	TOP			 	= 4'b0001,
				DOWN				= 4'b0010,
				UP		 			= 4'b0100,
				STOP				= 4'b1000;

localparam	FLAP_1 			= 2'd0,
				FLAP_2			= 2'd1,
				FLAP_3 			= 2'd2;
				
				
localparam TIME_START      =    20000;  // starting time to load when beginning to flap up
localparam TIME_STEP       =     5000;  // value to decrement or incremnt start time until above or below MAX or TERMINAL
localparam TIME_MAX        =   400000;  // start time for fall, end time for rise
localparam TIME_TERMINAL   =   150000;  // terminal time reached when falling down

reg [3:0] motion_state, prev_state;
reg [31:0] flap_elapsed, flap_start;

always @(posedge clk or posedge rst)
begin
	if (rst) begin
		motion_state 	<= DOWN;
		prev_state	 	<= DOWN;
		flap_elapsed 	<= TIME_MAX;
		flap_start		<= TIME_MAX;
		bird_state 		<= FLAP_1;
		birdY 			<= (480 - BIRD_SIZE_Y)/2;
	end else begin
		case (motion_state)
		
			TOP: begin
				prev_state 		<= TOP;
				
				flap_elapsed 	<= TIME_MAX;
				flap_start 		<= TIME_MAX;
				
				if (game_state != START_SCREEN || game_state != IN_GAME) begin
					motion_state <= STOP;
				end
				
				motion_state 	<= DOWN;
			end
			
			DOWN: begin
				prev_state	 	<= DOWN;
				bird_state 		<= FLAP_1;
				
				if (game_state != START_SCREEN || game_state != IN_GAME) begin
					motion_state <= STOP;
				end
				
				flap_elapsed 	<= flap_elapsed - 1;
				
				if (flap_elapsed == 0) begin					
					if (flap_start > TIME_TERMINAL) begin
						flap_start 		<= flap_start - TIME_STEP;
						flap_elapsed 	<= flap_start;
					end else begin
						flap_elapsed 	<= TIME_TERMINAL;
					end
					
					birdY <= birdY + 1;
				end
				
				if (flap || (game_state == START_SCREEN && birdY > 250)) begin
					motion_state 	<= UP;
					flap_start 		<= TIME_START;
					flap_elapsed 	<= TIME_START;
				end
			end
			
			UP: begin
				prev_state 		<= UP;
				
				if (flap_start <= (TIME_MAX/5) * 4)
					bird_state 	<= FLAP_3;
				else
					bird_state 	<= FLAP_2;
				
				if (game_state != START_SCREEN || game_state != IN_GAME) begin
					motion_state <= STOP;
				end
				
				flap_elapsed <= flap_elapsed - 1;
				
				if (flap_elapsed == 0) begin					
					if (flap_start <= TIME_MAX) begin
						flap_start 		<= flap_start + TIME_STEP;
						flap_elapsed 	<= flap_start;
						birdY 			<= birdY - 1;
					end else begin
						motion_state <= TOP;
					end
				end				
			end
			
			STOP: begin
				birdY <= birdY;
				if (game_state == START_SCREEN || game_state == IN_GAME) begin
					motion_state <= prev_state;
				end
			end
			
			default:	birdY <= birdY;
			
		endcase
	end
end

endmodule
		