module sprite_bitmap
(
	input [15:0] yofs, xofs,
	output [23:0] bit
);

reg [24*8 -1:0] bitarray [16:0];

assign bit = bitarray[yofs][xofs*24];

initial begin
	bitarray[0] 	= {24'hFFFFFF, 24'hFFFFFF, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[1] 	= {24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF, 24'hFF00FF, 24'hFF00FF, 24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[2] 	= {24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF, 24'hFF00FF, 24'hFF00FF, 24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[3] 	= {24'hFFFFFF, 24'hFFFFFF, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[4]		= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[5] 	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[6] 	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[7] 	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[8] 	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[9] 	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[10]	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[11]	= {24'h000000, 24'h000000, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'h000000, 24'h000000};
	bitarray[12]	= {24'hFFFFFF, 24'hFFFFFF, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[13]	= {24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF, 24'hFF00FF, 24'hFF00FF, 24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[14]	= {24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF, 24'hFF00FF, 24'hFF00FF, 24'hFFFFFF, 24'hFFFFFF, 24'hFFFFFF};
	bitarray[15]	= {24'hFFFFFF, 24'hFFFFFF, 24'h000000, 24'hFF00FF, 24'hFF00FF, 24'h000000, 24'hFFFFFF, 24'hFFFFFF};
end

endmodule
