module medals_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [4:0] col,
		output reg [23:0] colour_data
	);

	(* romstyle = "M4K" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: colour_data = 24'b111111110000000010010110;
		12'b000000000001: colour_data = 24'b111111110000000010010110;
		12'b000000000010: colour_data = 24'b111111110000000010010110;
		12'b000000000011: colour_data = 24'b111111110000000010010110;
		12'b000000000100: colour_data = 24'b111111110000000010010110;
		12'b000000000101: colour_data = 24'b111111110000000010010110;
		12'b000000000110: colour_data = 24'b111111110000000010010110;
		12'b000000000111: colour_data = 24'b111111110000000010010110;
		12'b000000001000: colour_data = 24'b101111011010001001000111;
		12'b000000001001: colour_data = 24'b101111011010001001000111;
		12'b000000001010: colour_data = 24'b101111011010001001000111;
		12'b000000001011: colour_data = 24'b101111011010001001000111;
		12'b000000001100: colour_data = 24'b101111011010001001000111;
		12'b000000001101: colour_data = 24'b101111011010001001000111;
		12'b000000001110: colour_data = 24'b111111110000000010010110;
		12'b000000001111: colour_data = 24'b111111110000000010010110;
		12'b000000010000: colour_data = 24'b111111110000000010010110;
		12'b000000010001: colour_data = 24'b111111110000000010010110;
		12'b000000010010: colour_data = 24'b111111110000000010010110;
		12'b000000010011: colour_data = 24'b111111110000000010010110;
		12'b000000010100: colour_data = 24'b111111110000000010010110;
		12'b000000010101: colour_data = 24'b111111110000000010010110;

		12'b000000100000: colour_data = 24'b111111110000000010010110;
		12'b000000100001: colour_data = 24'b111111110000000010010110;
		12'b000000100010: colour_data = 24'b111111110000000010010110;
		12'b000000100011: colour_data = 24'b111111110000000010010110;
		12'b000000100100: colour_data = 24'b111111110000000010010110;
		12'b000000100101: colour_data = 24'b111111110000000010010110;
		12'b000000100110: colour_data = 24'b101111011010001001000111;
		12'b000000100111: colour_data = 24'b101111011010001001000111;
		12'b000000101000: colour_data = 24'b111111111111111111111111;
		12'b000000101001: colour_data = 24'b111111111111111111111111;
		12'b000000101010: colour_data = 24'b111111111111111111111111;
		12'b000000101011: colour_data = 24'b111111111111111111111111;
		12'b000000101100: colour_data = 24'b111111111111111111111111;
		12'b000000101101: colour_data = 24'b111111111111111111111111;
		12'b000000101110: colour_data = 24'b101111011010001001000111;
		12'b000000101111: colour_data = 24'b101111011010001001000111;
		12'b000000110000: colour_data = 24'b111111110000000010010110;
		12'b000000110001: colour_data = 24'b111111110000000010010110;
		12'b000000110010: colour_data = 24'b111111110000000010010110;
		12'b000000110011: colour_data = 24'b111111110000000010010110;
		12'b000000110100: colour_data = 24'b111111110000000010010110;
		12'b000000110101: colour_data = 24'b111111110000000010010110;

		12'b000001000000: colour_data = 24'b111111110000000010010110;
		12'b000001000001: colour_data = 24'b111111110000000010010110;
		12'b000001000010: colour_data = 24'b111111110000000010010110;
		12'b000001000011: colour_data = 24'b111111110000000010010110;
		12'b000001000100: colour_data = 24'b101111011010001001000111;
		12'b000001000101: colour_data = 24'b101111011010001001000111;
		12'b000001000110: colour_data = 24'b111111111111111111111111;
		12'b000001000111: colour_data = 24'b111111111111111111111111;
		12'b000001001000: colour_data = 24'b111011011111001001100000;
		12'b000001001001: colour_data = 24'b111011011111001001100000;
		12'b000001001010: colour_data = 24'b111011011111001001100000;
		12'b000001001011: colour_data = 24'b111011011111001001100000;
		12'b000001001100: colour_data = 24'b111011011111001001100000;
		12'b000001001101: colour_data = 24'b111011011111001001100000;
		12'b000001001110: colour_data = 24'b111111111111111111111111;
		12'b000001001111: colour_data = 24'b111111111111111111111111;
		12'b000001010000: colour_data = 24'b101111011010001001000111;
		12'b000001010001: colour_data = 24'b101111011010001001000111;
		12'b000001010010: colour_data = 24'b111111110000000010010110;
		12'b000001010011: colour_data = 24'b111111110000000010010110;
		12'b000001010100: colour_data = 24'b111111110000000010010110;
		12'b000001010101: colour_data = 24'b111111110000000010010110;

		12'b000001100000: colour_data = 24'b111111110000000010010110;
		12'b000001100001: colour_data = 24'b111111110000000010010110;
		12'b000001100010: colour_data = 24'b111111110000000010010110;
		12'b000001100011: colour_data = 24'b101111011010001001000111;
		12'b000001100100: colour_data = 24'b111111111111111111111111;
		12'b000001100101: colour_data = 24'b111111111111111111111111;
		12'b000001100110: colour_data = 24'b111011011111001001100000;
		12'b000001100111: colour_data = 24'b111011011111001001100000;
		12'b000001101000: colour_data = 24'b111011011111001001100000;
		12'b000001101001: colour_data = 24'b111011011111001001100000;
		12'b000001101010: colour_data = 24'b111011011111001001100000;
		12'b000001101011: colour_data = 24'b111011011111001001100000;
		12'b000001101100: colour_data = 24'b111011011111001001100000;
		12'b000001101101: colour_data = 24'b111011011111001001100000;
		12'b000001101110: colour_data = 24'b111011011111001001100000;
		12'b000001101111: colour_data = 24'b111011011111001001100000;
		12'b000001110000: colour_data = 24'b111111111111111111111111;
		12'b000001110001: colour_data = 24'b111111111111111111111111;
		12'b000001110010: colour_data = 24'b101111011010001001000111;
		12'b000001110011: colour_data = 24'b111111110000000010010110;
		12'b000001110100: colour_data = 24'b111111110000000010010110;
		12'b000001110101: colour_data = 24'b111111110000000010010110;

		12'b000010000000: colour_data = 24'b111111110000000010010110;
		12'b000010000001: colour_data = 24'b111111110000000010010110;
		12'b000010000010: colour_data = 24'b101111011010001001000111;
		12'b000010000011: colour_data = 24'b111111111111111111111111;
		12'b000010000100: colour_data = 24'b111011011111001001100000;
		12'b000010000101: colour_data = 24'b111011011111001001100000;
		12'b000010000110: colour_data = 24'b111011011111001001100000;
		12'b000010000111: colour_data = 24'b111011011111001001100000;
		12'b000010001000: colour_data = 24'b111011011111001001100000;
		12'b000010001001: colour_data = 24'b111111111101101101011111;
		12'b000010001010: colour_data = 24'b111111111101101101011111;
		12'b000010001011: colour_data = 24'b111111111101101101011111;
		12'b000010001100: colour_data = 24'b111111111101101101011111;
		12'b000010001101: colour_data = 24'b111111111101101101011111;
		12'b000010001110: colour_data = 24'b111111111101101101011111;
		12'b000010001111: colour_data = 24'b111011011111001001100000;
		12'b000010010000: colour_data = 24'b111011011111001001100000;
		12'b000010010001: colour_data = 24'b111011011111001001100000;
		12'b000010010010: colour_data = 24'b111111111111111111111111;
		12'b000010010011: colour_data = 24'b101111011010001001000111;
		12'b000010010100: colour_data = 24'b111111110000000010010110;
		12'b000010010101: colour_data = 24'b111111110000000010010110;

		12'b000010100000: colour_data = 24'b111111110000000010010110;
		12'b000010100001: colour_data = 24'b111111110000000010010110;
		12'b000010100010: colour_data = 24'b101111011010001001000111;
		12'b000010100011: colour_data = 24'b111011011111001001100000;
		12'b000010100100: colour_data = 24'b111011011111001001100000;
		12'b000010100101: colour_data = 24'b111011011111001001100000;
		12'b000010100110: colour_data = 24'b111011011111001001100000;
		12'b000010100111: colour_data = 24'b111111111101101101011111;
		12'b000010101000: colour_data = 24'b111111111101101101011111;
		12'b000010101001: colour_data = 24'b111000111100001101010100;
		12'b000010101010: colour_data = 24'b111000111100001101010100;
		12'b000010101011: colour_data = 24'b111000111100001101010100;
		12'b000010101100: colour_data = 24'b111000111100001101010100;
		12'b000010101101: colour_data = 24'b111000111100001101010100;
		12'b000010101110: colour_data = 24'b111000111100001101010100;
		12'b000010101111: colour_data = 24'b111111111101101101011111;
		12'b000010110000: colour_data = 24'b111011011111001001100000;
		12'b000010110001: colour_data = 24'b111011011111001001100000;
		12'b000010110010: colour_data = 24'b111011011111001001100000;
		12'b000010110011: colour_data = 24'b101111011010001001000111;
		12'b000010110100: colour_data = 24'b111111110000000010010110;
		12'b000010110101: colour_data = 24'b111111110000000010010110;

		12'b000011000000: colour_data = 24'b111111110000000010010110;
		12'b000011000001: colour_data = 24'b101111011010001001000111;
		12'b000011000010: colour_data = 24'b111111111111111111111111;
		12'b000011000011: colour_data = 24'b111011011111001001100000;
		12'b000011000100: colour_data = 24'b111011011111001001100000;
		12'b000011000101: colour_data = 24'b111011011111001001100000;
		12'b000011000110: colour_data = 24'b111111111101101101011111;
		12'b000011000111: colour_data = 24'b111000111100001101010100;
		12'b000011001000: colour_data = 24'b111000111100001101010100;
		12'b000011001001: colour_data = 24'b111111111111111111111111;
		12'b000011001010: colour_data = 24'b111111111111111111111111;
		12'b000011001011: colour_data = 24'b111111111111111111111111;
		12'b000011001100: colour_data = 24'b111000111100001101010100;
		12'b000011001101: colour_data = 24'b111011011111001001100000;
		12'b000011001110: colour_data = 24'b111011011111001001100000;
		12'b000011001111: colour_data = 24'b111000111100001101010100;
		12'b000011010000: colour_data = 24'b111111111101101101011111;
		12'b000011010001: colour_data = 24'b111011011111001001100000;
		12'b000011010010: colour_data = 24'b111011011111001001100000;
		12'b000011010011: colour_data = 24'b111111111111111111111111;
		12'b000011010100: colour_data = 24'b101111011010001001000111;
		12'b000011010101: colour_data = 24'b111111110000000010010110;

		12'b000011100000: colour_data = 24'b111111110000000010010110;
		12'b000011100001: colour_data = 24'b101111011010001001000111;
		12'b000011100010: colour_data = 24'b111011011111001001100000;
		12'b000011100011: colour_data = 24'b111011011111001001100000;
		12'b000011100100: colour_data = 24'b111011011111001001100000;
		12'b000011100101: colour_data = 24'b111111111101101101011111;
		12'b000011100110: colour_data = 24'b111000111100001101010100;
		12'b000011100111: colour_data = 24'b111111111111111111111111;
		12'b000011101000: colour_data = 24'b111111111111111111111111;
		12'b000011101001: colour_data = 24'b111011011111001001100000;
		12'b000011101010: colour_data = 24'b111011011111001001100000;
		12'b000011101011: colour_data = 24'b111000111100001101010100;
		12'b000011101100: colour_data = 24'b111011011111001001100000;
		12'b000011101101: colour_data = 24'b111011011111001001100000;
		12'b000011101110: colour_data = 24'b111011011111001001100000;
		12'b000011101111: colour_data = 24'b111011011111001001100000;
		12'b000011110000: colour_data = 24'b111000111100001101010100;
		12'b000011110001: colour_data = 24'b111111111101101101011111;
		12'b000011110010: colour_data = 24'b111011011111001001100000;
		12'b000011110011: colour_data = 24'b111011011111001001100000;
		12'b000011110100: colour_data = 24'b101111011010001001000111;
		12'b000011110101: colour_data = 24'b111111110000000010010110;

		12'b000100000000: colour_data = 24'b101111011010001001000111;
		12'b000100000001: colour_data = 24'b111111111111111111111111;
		12'b000100000010: colour_data = 24'b111011011111001001100000;
		12'b000100000011: colour_data = 24'b111011011111001001100000;
		12'b000100000100: colour_data = 24'b111011011111001001100000;
		12'b000100000101: colour_data = 24'b111000111100001101010100;
		12'b000100000110: colour_data = 24'b111111111111111111111111;
		12'b000100000111: colour_data = 24'b111011011111001001100000;
		12'b000100001000: colour_data = 24'b111011011111001001100000;
		12'b000100001001: colour_data = 24'b111011011111001001100000;
		12'b000100001010: colour_data = 24'b111011011111001001100000;
		12'b000100001011: colour_data = 24'b111000111100001101010100;
		12'b000100001100: colour_data = 24'b111111111101101101011111;
		12'b000100001101: colour_data = 24'b111011011111001001100000;
		12'b000100001110: colour_data = 24'b111011011111001001100000;
		12'b000100001111: colour_data = 24'b111000111100001101010100;
		12'b000100010000: colour_data = 24'b111011011111001001100000;
		12'b000100010001: colour_data = 24'b111000111100001101010100;
		12'b000100010010: colour_data = 24'b111011011111001001100000;
		12'b000100010011: colour_data = 24'b111011011111001001100000;
		12'b000100010100: colour_data = 24'b111111111111111111111111;
		12'b000100010101: colour_data = 24'b101111011010001001000111;

		12'b000100100000: colour_data = 24'b101111011010001001000111;
		12'b000100100001: colour_data = 24'b111011011111001001100000;
		12'b000100100010: colour_data = 24'b111011011111001001100000;
		12'b000100100011: colour_data = 24'b111011011111001001100000;
		12'b000100100100: colour_data = 24'b111000111100001101010100;
		12'b000100100101: colour_data = 24'b111111111111111111111111;
		12'b000100100110: colour_data = 24'b111011011111001001100000;
		12'b000100100111: colour_data = 24'b111011011111001001100000;
		12'b000100101000: colour_data = 24'b111011011111001001100000;
		12'b000100101001: colour_data = 24'b111011011111001001100000;
		12'b000100101010: colour_data = 24'b111011011111001001100000;
		12'b000100101011: colour_data = 24'b111000111100001101010100;
		12'b000100101100: colour_data = 24'b111111111101101101011111;
		12'b000100101101: colour_data = 24'b111011011111001001100000;
		12'b000100101110: colour_data = 24'b111011011111001001100000;
		12'b000100101111: colour_data = 24'b111000111100001101010100;
		12'b000100110000: colour_data = 24'b111011011111001001100000;
		12'b000100110001: colour_data = 24'b111000111100001101010100;
		12'b000100110010: colour_data = 24'b111011011111001001100000;
		12'b000100110011: colour_data = 24'b111011011111001001100000;
		12'b000100110100: colour_data = 24'b111011011111001001100000;
		12'b000100110101: colour_data = 24'b101111011010001001000111;

		12'b000101000000: colour_data = 24'b101111011010001001000111;
		12'b000101000001: colour_data = 24'b111011011111001001100000;
		12'b000101000010: colour_data = 24'b111011011111001001100000;
		12'b000101000011: colour_data = 24'b111011011111001001100000;
		12'b000101000100: colour_data = 24'b111000111100001101010100;
		12'b000101000101: colour_data = 24'b111011011111001001100000;
		12'b000101000110: colour_data = 24'b111011011111001001100000;
		12'b000101000111: colour_data = 24'b111011011111001001100000;
		12'b000101001000: colour_data = 24'b111011011111001001100000;
		12'b000101001001: colour_data = 24'b111011011111001001100000;
		12'b000101001010: colour_data = 24'b111011011111001001100000;
		12'b000101001011: colour_data = 24'b111011011111001001100000;
		12'b000101001100: colour_data = 24'b111000111100001101010100;
		12'b000101001101: colour_data = 24'b111111111101101101011111;
		12'b000101001110: colour_data = 24'b111011011111001001100000;
		12'b000101001111: colour_data = 24'b111011011111001001100000;
		12'b000101010000: colour_data = 24'b111011011111001001100000;
		12'b000101010001: colour_data = 24'b111000111100001101010100;
		12'b000101010010: colour_data = 24'b111111111101101101011111;
		12'b000101010011: colour_data = 24'b111011011111001001100000;
		12'b000101010100: colour_data = 24'b111011011111001001100000;
		12'b000101010101: colour_data = 24'b101111011010001001000111;

		12'b000101100000: colour_data = 24'b101111011010001001000111;
		12'b000101100001: colour_data = 24'b111011011111001001100000;
		12'b000101100010: colour_data = 24'b111011011111001001100000;
		12'b000101100011: colour_data = 24'b111111111101101101011111;
		12'b000101100100: colour_data = 24'b111000111100001101010100;
		12'b000101100101: colour_data = 24'b111000111100001101010100;
		12'b000101100110: colour_data = 24'b111000111100001101010100;
		12'b000101100111: colour_data = 24'b111000111100001101010100;
		12'b000101101000: colour_data = 24'b111000111100001101010100;
		12'b000101101001: colour_data = 24'b111011011111001001100000;
		12'b000101101010: colour_data = 24'b111011011111001001100000;
		12'b000101101011: colour_data = 24'b111011011111001001100000;
		12'b000101101100: colour_data = 24'b111011011111001001100000;
		12'b000101101101: colour_data = 24'b111000111100001101010100;
		12'b000101101110: colour_data = 24'b111000111100001101010100;
		12'b000101101111: colour_data = 24'b111000111100001101010100;
		12'b000101110000: colour_data = 24'b111000111100001101010100;
		12'b000101110001: colour_data = 24'b111000111100001101010100;
		12'b000101110010: colour_data = 24'b111000111100001101010100;
		12'b000101110011: colour_data = 24'b111111111101101101011111;
		12'b000101110100: colour_data = 24'b111011011111001001100000;
		12'b000101110101: colour_data = 24'b101111011010001001000111;

		12'b000110000000: colour_data = 24'b101111011010001001000111;
		12'b000110000001: colour_data = 24'b111011011111001001100000;
		12'b000110000010: colour_data = 24'b111011011111001001100000;
		12'b000110000011: colour_data = 24'b111000111100001101010100;
		12'b000110000100: colour_data = 24'b111011011111001001100000;
		12'b000110000101: colour_data = 24'b111111111111111111111111;
		12'b000110000110: colour_data = 24'b111111111111111111111111;
		12'b000110000111: colour_data = 24'b111111111111111111111111;
		12'b000110001000: colour_data = 24'b111011011111001001100000;
		12'b000110001001: colour_data = 24'b111000111100001101010100;
		12'b000110001010: colour_data = 24'b111011011111001001100000;
		12'b000110001011: colour_data = 24'b111011011111001001100000;
		12'b000110001100: colour_data = 24'b111000111100001101010100;
		12'b000110001101: colour_data = 24'b111011011111001001100000;
		12'b000110001110: colour_data = 24'b111011011111001001100000;
		12'b000110001111: colour_data = 24'b111011011111001001100000;
		12'b000110010000: colour_data = 24'b111011011111001001100000;
		12'b000110010001: colour_data = 24'b111011011111001001100000;
		12'b000110010010: colour_data = 24'b111011011111001001100000;
		12'b000110010011: colour_data = 24'b111000111100001101010100;
		12'b000110010100: colour_data = 24'b111011011111001001100000;
		12'b000110010101: colour_data = 24'b101111011010001001000111;

		12'b000110100000: colour_data = 24'b101111011010001001000111;
		12'b000110100001: colour_data = 24'b111111111101101101011111;
		12'b000110100010: colour_data = 24'b111011011111001001100000;
		12'b000110100011: colour_data = 24'b111000111100001101010100;
		12'b000110100100: colour_data = 24'b111111111111111111111111;
		12'b000110100101: colour_data = 24'b111111111111111111111111;
		12'b000110100110: colour_data = 24'b111111111111111111111111;
		12'b000110100111: colour_data = 24'b111111111111111111111111;
		12'b000110101000: colour_data = 24'b111000111100001101010100;
		12'b000110101001: colour_data = 24'b111111111101101101011111;
		12'b000110101010: colour_data = 24'b111111111101101101011111;
		12'b000110101011: colour_data = 24'b111000111100001101010100;
		12'b000110101100: colour_data = 24'b111011011111001001100000;
		12'b000110101101: colour_data = 24'b111000111100001101010100;
		12'b000110101110: colour_data = 24'b111000111100001101010100;
		12'b000110101111: colour_data = 24'b111000111100001101010100;
		12'b000110110000: colour_data = 24'b111000111100001101010100;
		12'b000110110001: colour_data = 24'b111000111100001101010100;
		12'b000110110010: colour_data = 24'b111000111100001101010100;
		12'b000110110011: colour_data = 24'b111111111111111111111111;
		12'b000110110100: colour_data = 24'b111111111101101101011111;
		12'b000110110101: colour_data = 24'b101111011010001001000111;

		12'b000111000000: colour_data = 24'b111111110000000010010110;
		12'b000111000001: colour_data = 24'b101111011010001001000111;
		12'b000111000010: colour_data = 24'b111011011111001001100000;
		12'b000111000011: colour_data = 24'b111000111100001101010100;
		12'b000111000100: colour_data = 24'b111111111111111111111111;
		12'b000111000101: colour_data = 24'b111111111111111111111111;
		12'b000111000110: colour_data = 24'b111011011111001001100000;
		12'b000111000111: colour_data = 24'b111000111100001101010100;
		12'b000111001000: colour_data = 24'b111111111101101101011111;
		12'b000111001001: colour_data = 24'b111111111101101101011111;
		12'b000111001010: colour_data = 24'b111111111101101101011111;
		12'b000111001011: colour_data = 24'b111111111101101101011111;
		12'b000111001100: colour_data = 24'b111000111100001101010100;
		12'b000111001101: colour_data = 24'b111011011111001001100000;
		12'b000111001110: colour_data = 24'b111011011111001001100000;
		12'b000111001111: colour_data = 24'b111011011111001001100000;
		12'b000111010000: colour_data = 24'b111011011111001001100000;
		12'b000111010001: colour_data = 24'b111011011111001001100000;
		12'b000111010010: colour_data = 24'b111000111100001101010100;
		12'b000111010011: colour_data = 24'b111011011111001001100000;
		12'b000111010100: colour_data = 24'b101111011010001001000111;
		12'b000111010101: colour_data = 24'b111111110000000010010110;

		12'b000111100000: colour_data = 24'b111111110000000010010110;
		12'b000111100001: colour_data = 24'b101111011010001001000111;
		12'b000111100010: colour_data = 24'b111111111101101101011111;
		12'b000111100011: colour_data = 24'b111111111111111111111111;
		12'b000111100100: colour_data = 24'b111000111100001101010100;
		12'b000111100101: colour_data = 24'b111000111100001101010100;
		12'b000111100110: colour_data = 24'b111000111100001101010100;
		12'b000111100111: colour_data = 24'b111000111100001101010100;
		12'b000111101000: colour_data = 24'b111111111101101101011111;
		12'b000111101001: colour_data = 24'b111111111101101101011111;
		12'b000111101010: colour_data = 24'b111111111101101101011111;
		12'b000111101011: colour_data = 24'b111111111101101101011111;
		12'b000111101100: colour_data = 24'b111111111101101101011111;
		12'b000111101101: colour_data = 24'b111000111100001101010100;
		12'b000111101110: colour_data = 24'b111000111100001101010100;
		12'b000111101111: colour_data = 24'b111000111100001101010100;
		12'b000111110000: colour_data = 24'b111000111100001101010100;
		12'b000111110001: colour_data = 24'b111000111100001101010100;
		12'b000111110010: colour_data = 24'b111111111111111111111111;
		12'b000111110011: colour_data = 24'b111111111101101101011111;
		12'b000111110100: colour_data = 24'b101111011010001001000111;
		12'b000111110101: colour_data = 24'b111111110000000010010110;

		12'b001000000000: colour_data = 24'b111111110000000010010110;
		12'b001000000001: colour_data = 24'b111111110000000010010110;
		12'b001000000010: colour_data = 24'b101111011010001001000111;
		12'b001000000011: colour_data = 24'b111011011111001001100000;
		12'b001000000100: colour_data = 24'b111111111111111111111111;
		12'b001000000101: colour_data = 24'b111111111111111111111111;
		12'b001000000110: colour_data = 24'b111111111111111111111111;
		12'b001000000111: colour_data = 24'b111111111111111111111111;
		12'b001000001000: colour_data = 24'b111000111100001101010100;
		12'b001000001001: colour_data = 24'b111000111100001101010100;
		12'b001000001010: colour_data = 24'b111000111100001101010100;
		12'b001000001011: colour_data = 24'b111000111100001101010100;
		12'b001000001100: colour_data = 24'b111000111100001101010100;
		12'b001000001101: colour_data = 24'b111111111111111111111111;
		12'b001000001110: colour_data = 24'b111111111111111111111111;
		12'b001000001111: colour_data = 24'b111111111111111111111111;
		12'b001000010000: colour_data = 24'b111111111111111111111111;
		12'b001000010001: colour_data = 24'b111111111111111111111111;
		12'b001000010010: colour_data = 24'b111011011111001001100000;
		12'b001000010011: colour_data = 24'b101111011010001001000111;
		12'b001000010100: colour_data = 24'b111111110000000010010110;
		12'b001000010101: colour_data = 24'b111111110000000010010110;

		12'b001000100000: colour_data = 24'b111111110000000010010110;
		12'b001000100001: colour_data = 24'b111111110000000010010110;
		12'b001000100010: colour_data = 24'b101111011010001001000111;
		12'b001000100011: colour_data = 24'b111111111101101101011111;
		12'b001000100100: colour_data = 24'b111011011111001001100000;
		12'b001000100101: colour_data = 24'b111011011111001001100000;
		12'b001000100110: colour_data = 24'b111011011111001001100000;
		12'b001000100111: colour_data = 24'b111011011111001001100000;
		12'b001000101000: colour_data = 24'b111111111111111111111111;
		12'b001000101001: colour_data = 24'b111111111111111111111111;
		12'b001000101010: colour_data = 24'b111111111111111111111111;
		12'b001000101011: colour_data = 24'b111111111111111111111111;
		12'b001000101100: colour_data = 24'b111111111111111111111111;
		12'b001000101101: colour_data = 24'b111011011111001001100000;
		12'b001000101110: colour_data = 24'b111011011111001001100000;
		12'b001000101111: colour_data = 24'b111011011111001001100000;
		12'b001000110000: colour_data = 24'b111011011111001001100000;
		12'b001000110001: colour_data = 24'b111011011111001001100000;
		12'b001000110010: colour_data = 24'b111111111101101101011111;
		12'b001000110011: colour_data = 24'b101111011010001001000111;
		12'b001000110100: colour_data = 24'b111111110000000010010110;
		12'b001000110101: colour_data = 24'b111111110000000010010110;

		12'b001001000000: colour_data = 24'b111111110000000010010110;
		12'b001001000001: colour_data = 24'b111111110000000010010110;
		12'b001001000010: colour_data = 24'b111111110000000010010110;
		12'b001001000011: colour_data = 24'b101111011010001001000111;
		12'b001001000100: colour_data = 24'b111111111101101101011111;
		12'b001001000101: colour_data = 24'b111111111101101101011111;
		12'b001001000110: colour_data = 24'b111011011111001001100000;
		12'b001001000111: colour_data = 24'b111011011111001001100000;
		12'b001001001000: colour_data = 24'b111011011111001001100000;
		12'b001001001001: colour_data = 24'b111011011111001001100000;
		12'b001001001010: colour_data = 24'b111011011111001001100000;
		12'b001001001011: colour_data = 24'b111011011111001001100000;
		12'b001001001100: colour_data = 24'b111011011111001001100000;
		12'b001001001101: colour_data = 24'b111011011111001001100000;
		12'b001001001110: colour_data = 24'b111011011111001001100000;
		12'b001001001111: colour_data = 24'b111011011111001001100000;
		12'b001001010000: colour_data = 24'b111111111101101101011111;
		12'b001001010001: colour_data = 24'b111111111101101101011111;
		12'b001001010010: colour_data = 24'b101111011010001001000111;
		12'b001001010011: colour_data = 24'b111111110000000010010110;
		12'b001001010100: colour_data = 24'b111111110000000010010110;
		12'b001001010101: colour_data = 24'b111111110000000010010110;

		12'b001001100000: colour_data = 24'b111111110000000010010110;
		12'b001001100001: colour_data = 24'b111111110000000010010110;
		12'b001001100010: colour_data = 24'b111111110000000010010110;
		12'b001001100011: colour_data = 24'b111111110000000010010110;
		12'b001001100100: colour_data = 24'b101111011010001001000111;
		12'b001001100101: colour_data = 24'b101111011010001001000111;
		12'b001001100110: colour_data = 24'b111111111101101101011111;
		12'b001001100111: colour_data = 24'b111111111101101101011111;
		12'b001001101000: colour_data = 24'b111011011111001001100000;
		12'b001001101001: colour_data = 24'b111011011111001001100000;
		12'b001001101010: colour_data = 24'b111011011111001001100000;
		12'b001001101011: colour_data = 24'b111011011111001001100000;
		12'b001001101100: colour_data = 24'b111011011111001001100000;
		12'b001001101101: colour_data = 24'b111011011111001001100000;
		12'b001001101110: colour_data = 24'b111111111101101101011111;
		12'b001001101111: colour_data = 24'b111111111101101101011111;
		12'b001001110000: colour_data = 24'b101111011010001001000111;
		12'b001001110001: colour_data = 24'b101111011010001001000111;
		12'b001001110010: colour_data = 24'b111111110000000010010110;
		12'b001001110011: colour_data = 24'b111111110000000010010110;
		12'b001001110100: colour_data = 24'b111111110000000010010110;
		12'b001001110101: colour_data = 24'b111111110000000010010110;

		12'b001010000000: colour_data = 24'b111111110000000010010110;
		12'b001010000001: colour_data = 24'b111111110000000010010110;
		12'b001010000010: colour_data = 24'b111111110000000010010110;
		12'b001010000011: colour_data = 24'b111111110000000010010110;
		12'b001010000100: colour_data = 24'b111111110000000010010110;
		12'b001010000101: colour_data = 24'b111111110000000010010110;
		12'b001010000110: colour_data = 24'b101111011010001001000111;
		12'b001010000111: colour_data = 24'b101111011010001001000111;
		12'b001010001000: colour_data = 24'b111111111101101101011111;
		12'b001010001001: colour_data = 24'b111111111101101101011111;
		12'b001010001010: colour_data = 24'b111111111101101101011111;
		12'b001010001011: colour_data = 24'b111111111101101101011111;
		12'b001010001100: colour_data = 24'b111111111101101101011111;
		12'b001010001101: colour_data = 24'b111111111101101101011111;
		12'b001010001110: colour_data = 24'b101111011010001001000111;
		12'b001010001111: colour_data = 24'b101111011010001001000111;
		12'b001010010000: colour_data = 24'b111111110000000010010110;
		12'b001010010001: colour_data = 24'b111111110000000010010110;
		12'b001010010010: colour_data = 24'b111111110000000010010110;
		12'b001010010011: colour_data = 24'b111111110000000010010110;
		12'b001010010100: colour_data = 24'b111111110000000010010110;
		12'b001010010101: colour_data = 24'b111111110000000010010110;

		12'b001010100000: colour_data = 24'b111111110000000010010110;
		12'b001010100001: colour_data = 24'b111111110000000010010110;
		12'b001010100010: colour_data = 24'b111111110000000010010110;
		12'b001010100011: colour_data = 24'b111111110000000010010110;
		12'b001010100100: colour_data = 24'b111111110000000010010110;
		12'b001010100101: colour_data = 24'b111111110000000010010110;
		12'b001010100110: colour_data = 24'b111111110000000010010110;
		12'b001010100111: colour_data = 24'b111111110000000010010110;
		12'b001010101000: colour_data = 24'b101111011010001001000111;
		12'b001010101001: colour_data = 24'b101111011010001001000111;
		12'b001010101010: colour_data = 24'b101111011010001001000111;
		12'b001010101011: colour_data = 24'b101111011010001001000111;
		12'b001010101100: colour_data = 24'b101111011010001001000111;
		12'b001010101101: colour_data = 24'b101111011010001001000111;
		12'b001010101110: colour_data = 24'b111111110000000010010110;
		12'b001010101111: colour_data = 24'b111111110000000010010110;
		12'b001010110000: colour_data = 24'b111111110000000010010110;
		12'b001010110001: colour_data = 24'b111111110000000010010110;
		12'b001010110010: colour_data = 24'b111111110000000010010110;
		12'b001010110011: colour_data = 24'b111111110000000010010110;
		12'b001010110100: colour_data = 24'b111111110000000010010110;
		12'b001010110101: colour_data = 24'b111111110000000010010110;

		12'b001011000000: colour_data = 24'b111111110000000010010110;
		12'b001011000001: colour_data = 24'b111111110000000010010110;
		12'b001011000010: colour_data = 24'b111111110000000010010110;
		12'b001011000011: colour_data = 24'b111111110000000010010110;
		12'b001011000100: colour_data = 24'b111111110000000010010110;
		12'b001011000101: colour_data = 24'b111111110000000010010110;
		12'b001011000110: colour_data = 24'b111111110000000010010110;
		12'b001011000111: colour_data = 24'b111111110000000010010110;
		12'b001011001000: colour_data = 24'b100001000111111101111111;
		12'b001011001001: colour_data = 24'b100001000111111101111111;
		12'b001011001010: colour_data = 24'b100001000111111101111111;
		12'b001011001011: colour_data = 24'b100001000111111101111111;
		12'b001011001100: colour_data = 24'b100001000111111101111111;
		12'b001011001101: colour_data = 24'b100001000111111101111111;
		12'b001011001110: colour_data = 24'b111111110000000010010110;
		12'b001011001111: colour_data = 24'b111111110000000010010110;
		12'b001011010000: colour_data = 24'b111111110000000010010110;
		12'b001011010001: colour_data = 24'b111111110000000010010110;
		12'b001011010010: colour_data = 24'b111111110000000010010110;
		12'b001011010011: colour_data = 24'b111111110000000010010110;
		12'b001011010100: colour_data = 24'b111111110000000010010110;
		12'b001011010101: colour_data = 24'b111111110000000010010110;

		12'b001011100000: colour_data = 24'b111111110000000010010110;
		12'b001011100001: colour_data = 24'b111111110000000010010110;
		12'b001011100010: colour_data = 24'b111111110000000010010110;
		12'b001011100011: colour_data = 24'b111111110000000010010110;
		12'b001011100100: colour_data = 24'b111111110000000010010110;
		12'b001011100101: colour_data = 24'b111111110000000010010110;
		12'b001011100110: colour_data = 24'b100001000111111101111111;
		12'b001011100111: colour_data = 24'b100001000111111101111111;
		12'b001011101000: colour_data = 24'b111111111111111111111111;
		12'b001011101001: colour_data = 24'b111111111111111111111111;
		12'b001011101010: colour_data = 24'b111111111111111111111111;
		12'b001011101011: colour_data = 24'b111111111111111111111111;
		12'b001011101100: colour_data = 24'b111111111111111111111111;
		12'b001011101101: colour_data = 24'b111111111111111111111111;
		12'b001011101110: colour_data = 24'b100001000111111101111111;
		12'b001011101111: colour_data = 24'b100001000111111101111111;
		12'b001011110000: colour_data = 24'b111111110000000010010110;
		12'b001011110001: colour_data = 24'b111111110000000010010110;
		12'b001011110010: colour_data = 24'b111111110000000010010110;
		12'b001011110011: colour_data = 24'b111111110000000010010110;
		12'b001011110100: colour_data = 24'b111111110000000010010110;
		12'b001011110101: colour_data = 24'b111111110000000010010110;

		12'b001100000000: colour_data = 24'b111111110000000010010110;
		12'b001100000001: colour_data = 24'b111111110000000010010110;
		12'b001100000010: colour_data = 24'b111111110000000010010110;
		12'b001100000011: colour_data = 24'b111111110000000010010110;
		12'b001100000100: colour_data = 24'b100001000111111101111111;
		12'b001100000101: colour_data = 24'b100001000111111101111111;
		12'b001100000110: colour_data = 24'b111111111111111111111111;
		12'b001100000111: colour_data = 24'b111111111111111111111111;
		12'b001100001000: colour_data = 24'b111010011110000111100001;
		12'b001100001001: colour_data = 24'b111010011110000111100001;
		12'b001100001010: colour_data = 24'b111010011110000111100001;
		12'b001100001011: colour_data = 24'b111010011110000111100001;
		12'b001100001100: colour_data = 24'b111010011110000111100001;
		12'b001100001101: colour_data = 24'b111010011110000111100001;
		12'b001100001110: colour_data = 24'b111111111111111111111111;
		12'b001100001111: colour_data = 24'b111111111111111111111111;
		12'b001100010000: colour_data = 24'b100001000111111101111111;
		12'b001100010001: colour_data = 24'b100001000111111101111111;
		12'b001100010010: colour_data = 24'b111111110000000010010110;
		12'b001100010011: colour_data = 24'b111111110000000010010110;
		12'b001100010100: colour_data = 24'b111111110000000010010110;
		12'b001100010101: colour_data = 24'b111111110000000010010110;

		12'b001100100000: colour_data = 24'b111111110000000010010110;
		12'b001100100001: colour_data = 24'b111111110000000010010110;
		12'b001100100010: colour_data = 24'b111111110000000010010110;
		12'b001100100011: colour_data = 24'b100001000111111101111111;
		12'b001100100100: colour_data = 24'b111111111111111111111111;
		12'b001100100101: colour_data = 24'b111111111111111111111111;
		12'b001100100110: colour_data = 24'b111010011110000111100001;
		12'b001100100111: colour_data = 24'b111010011110000111100001;
		12'b001100101000: colour_data = 24'b111010011110000111100001;
		12'b001100101001: colour_data = 24'b111010011110000111100001;
		12'b001100101010: colour_data = 24'b111010011110000111100001;
		12'b001100101011: colour_data = 24'b111010011110000111100001;
		12'b001100101100: colour_data = 24'b111010011110000111100001;
		12'b001100101101: colour_data = 24'b111010011110000111100001;
		12'b001100101110: colour_data = 24'b111010011110000111100001;
		12'b001100101111: colour_data = 24'b111010011110000111100001;
		12'b001100110000: colour_data = 24'b111111111111111111111111;
		12'b001100110001: colour_data = 24'b111111111111111111111111;
		12'b001100110010: colour_data = 24'b100001000111111101111111;
		12'b001100110011: colour_data = 24'b111111110000000010010110;
		12'b001100110100: colour_data = 24'b111111110000000010010110;
		12'b001100110101: colour_data = 24'b111111110000000010010110;

		12'b001101000000: colour_data = 24'b111111110000000010010110;
		12'b001101000001: colour_data = 24'b111111110000000010010110;
		12'b001101000010: colour_data = 24'b100001000111111101111111;
		12'b001101000011: colour_data = 24'b111111111111111111111111;
		12'b001101000100: colour_data = 24'b111010011110000111100001;
		12'b001101000101: colour_data = 24'b111010011110000111100001;
		12'b001101000110: colour_data = 24'b111010011110000111100001;
		12'b001101000111: colour_data = 24'b111010011110000111100001;
		12'b001101001000: colour_data = 24'b111010011110000111100001;
		12'b001101001001: colour_data = 24'b110010001100000011000000;
		12'b001101001010: colour_data = 24'b110010001100000011000000;
		12'b001101001011: colour_data = 24'b110010001100000011000000;
		12'b001101001100: colour_data = 24'b110010001100000011000000;
		12'b001101001101: colour_data = 24'b110010001100000011000000;
		12'b001101001110: colour_data = 24'b110010001100000011000000;
		12'b001101001111: colour_data = 24'b111010011110000111100001;
		12'b001101010000: colour_data = 24'b111010011110000111100001;
		12'b001101010001: colour_data = 24'b111010011110000111100001;
		12'b001101010010: colour_data = 24'b111111111111111111111111;
		12'b001101010011: colour_data = 24'b100001000111111101111111;
		12'b001101010100: colour_data = 24'b111111110000000010010110;
		12'b001101010101: colour_data = 24'b111111110000000010010110;

		12'b001101100000: colour_data = 24'b111111110000000010010110;
		12'b001101100001: colour_data = 24'b111111110000000010010110;
		12'b001101100010: colour_data = 24'b100001000111111101111111;
		12'b001101100011: colour_data = 24'b111010011110000111100001;
		12'b001101100100: colour_data = 24'b111010011110000111100001;
		12'b001101100101: colour_data = 24'b111010011110000111100001;
		12'b001101100110: colour_data = 24'b111010011110000111100001;
		12'b001101100111: colour_data = 24'b110010001100000011000000;
		12'b001101101000: colour_data = 24'b110010001100000011000000;
		12'b001101101001: colour_data = 24'b100111011001100010011000;
		12'b001101101010: colour_data = 24'b100111011001100010011000;
		12'b001101101011: colour_data = 24'b100111011001100010011000;
		12'b001101101100: colour_data = 24'b100111011001100010011000;
		12'b001101101101: colour_data = 24'b100111011001100010011000;
		12'b001101101110: colour_data = 24'b100111011001100010011000;
		12'b001101101111: colour_data = 24'b110010001100000011000000;
		12'b001101110000: colour_data = 24'b111010011110000111100001;
		12'b001101110001: colour_data = 24'b111010011110000111100001;
		12'b001101110010: colour_data = 24'b111010011110000111100001;
		12'b001101110011: colour_data = 24'b100001000111111101111111;
		12'b001101110100: colour_data = 24'b111111110000000010010110;
		12'b001101110101: colour_data = 24'b111111110000000010010110;

		12'b001110000000: colour_data = 24'b111111110000000010010110;
		12'b001110000001: colour_data = 24'b100001000111111101111111;
		12'b001110000010: colour_data = 24'b111111111111111111111111;
		12'b001110000011: colour_data = 24'b111010011110000111100001;
		12'b001110000100: colour_data = 24'b111010011110000111100001;
		12'b001110000101: colour_data = 24'b111010011110000111100001;
		12'b001110000110: colour_data = 24'b110010001100000011000000;
		12'b001110000111: colour_data = 24'b100111011001100010011000;
		12'b001110001000: colour_data = 24'b100111011001100010011000;
		12'b001110001001: colour_data = 24'b111111111111111111111111;
		12'b001110001010: colour_data = 24'b111111111111111111111111;
		12'b001110001011: colour_data = 24'b111111111111111111111111;
		12'b001110001100: colour_data = 24'b100111011001100010011000;
		12'b001110001101: colour_data = 24'b111010011110000111100001;
		12'b001110001110: colour_data = 24'b111010011110000111100001;
		12'b001110001111: colour_data = 24'b100111011001100010011000;
		12'b001110010000: colour_data = 24'b110010001100000011000000;
		12'b001110010001: colour_data = 24'b111010011110000111100001;
		12'b001110010010: colour_data = 24'b111010011110000111100001;
		12'b001110010011: colour_data = 24'b111111111111111111111111;
		12'b001110010100: colour_data = 24'b100001000111111101111111;
		12'b001110010101: colour_data = 24'b111111110000000010010110;

		12'b001110100000: colour_data = 24'b111111110000000010010110;
		12'b001110100001: colour_data = 24'b100001000111111101111111;
		12'b001110100010: colour_data = 24'b111010011110000111100001;
		12'b001110100011: colour_data = 24'b111010011110000111100001;
		12'b001110100100: colour_data = 24'b111010011110000111100001;
		12'b001110100101: colour_data = 24'b110010001100000011000000;
		12'b001110100110: colour_data = 24'b100111011001100010011000;
		12'b001110100111: colour_data = 24'b111111111111111111111111;
		12'b001110101000: colour_data = 24'b111111111111111111111111;
		12'b001110101001: colour_data = 24'b111010011110000111100001;
		12'b001110101010: colour_data = 24'b111010011110000111100001;
		12'b001110101011: colour_data = 24'b100111011001100010011000;
		12'b001110101100: colour_data = 24'b111010011110000111100001;
		12'b001110101101: colour_data = 24'b111010011110000111100001;
		12'b001110101110: colour_data = 24'b111010011110000111100001;
		12'b001110101111: colour_data = 24'b111010011110000111100001;
		12'b001110110000: colour_data = 24'b100111011001100010011000;
		12'b001110110001: colour_data = 24'b110010001100000011000000;
		12'b001110110010: colour_data = 24'b111010011110000111100001;
		12'b001110110011: colour_data = 24'b111010011110000111100001;
		12'b001110110100: colour_data = 24'b100001000111111101111111;
		12'b001110110101: colour_data = 24'b111111110000000010010110;

		12'b001111000000: colour_data = 24'b100001000111111101111111;
		12'b001111000001: colour_data = 24'b111111111111111111111111;
		12'b001111000010: colour_data = 24'b111010011110000111100001;
		12'b001111000011: colour_data = 24'b111010011110000111100001;
		12'b001111000100: colour_data = 24'b111010011110000111100001;
		12'b001111000101: colour_data = 24'b100111011001100010011000;
		12'b001111000110: colour_data = 24'b111111111111111111111111;
		12'b001111000111: colour_data = 24'b111010011110000111100001;
		12'b001111001000: colour_data = 24'b111010011110000111100001;
		12'b001111001001: colour_data = 24'b111010011110000111100001;
		12'b001111001010: colour_data = 24'b111010011110000111100001;
		12'b001111001011: colour_data = 24'b100111011001100010011000;
		12'b001111001100: colour_data = 24'b110010001100000011000000;
		12'b001111001101: colour_data = 24'b111010011110000111100001;
		12'b001111001110: colour_data = 24'b111010011110000111100001;
		12'b001111001111: colour_data = 24'b100111011001100010011000;
		12'b001111010000: colour_data = 24'b111010011110000111100001;
		12'b001111010001: colour_data = 24'b100111011001100010011000;
		12'b001111010010: colour_data = 24'b111010011110000111100001;
		12'b001111010011: colour_data = 24'b111010011110000111100001;
		12'b001111010100: colour_data = 24'b111111111111111111111111;
		12'b001111010101: colour_data = 24'b100001000111111101111111;

		12'b001111100000: colour_data = 24'b100001000111111101111111;
		12'b001111100001: colour_data = 24'b111010011110000111100001;
		12'b001111100010: colour_data = 24'b111010011110000111100001;
		12'b001111100011: colour_data = 24'b111010011110000111100001;
		12'b001111100100: colour_data = 24'b100111011001100010011000;
		12'b001111100101: colour_data = 24'b111111111111111111111111;
		12'b001111100110: colour_data = 24'b111010011110000111100001;
		12'b001111100111: colour_data = 24'b111010011110000111100001;
		12'b001111101000: colour_data = 24'b111010011110000111100001;
		12'b001111101001: colour_data = 24'b111010011110000111100001;
		12'b001111101010: colour_data = 24'b111010011110000111100001;
		12'b001111101011: colour_data = 24'b100111011001100010011000;
		12'b001111101100: colour_data = 24'b110010001100000011000000;
		12'b001111101101: colour_data = 24'b111010011110000111100001;
		12'b001111101110: colour_data = 24'b111010011110000111100001;
		12'b001111101111: colour_data = 24'b100111011001100010011000;
		12'b001111110000: colour_data = 24'b111010011110000111100001;
		12'b001111110001: colour_data = 24'b100111011001100010011000;
		12'b001111110010: colour_data = 24'b111010011110000111100001;
		12'b001111110011: colour_data = 24'b111010011110000111100001;
		12'b001111110100: colour_data = 24'b111010011110000111100001;
		12'b001111110101: colour_data = 24'b100001000111111101111111;

		12'b010000000000: colour_data = 24'b100001000111111101111111;
		12'b010000000001: colour_data = 24'b111010011110000111100001;
		12'b010000000010: colour_data = 24'b111010011110000111100001;
		12'b010000000011: colour_data = 24'b111010011110000111100001;
		12'b010000000100: colour_data = 24'b100111011001100010011000;
		12'b010000000101: colour_data = 24'b111010011110000111100001;
		12'b010000000110: colour_data = 24'b111010011110000111100001;
		12'b010000000111: colour_data = 24'b111010011110000111100001;
		12'b010000001000: colour_data = 24'b111010011110000111100001;
		12'b010000001001: colour_data = 24'b111010011110000111100001;
		12'b010000001010: colour_data = 24'b111010011110000111100001;
		12'b010000001011: colour_data = 24'b111010011110000111100001;
		12'b010000001100: colour_data = 24'b100111011001100010011000;
		12'b010000001101: colour_data = 24'b110010001100000011000000;
		12'b010000001110: colour_data = 24'b111010011110000111100001;
		12'b010000001111: colour_data = 24'b111010011110000111100001;
		12'b010000010000: colour_data = 24'b111010011110000111100001;
		12'b010000010001: colour_data = 24'b100111011001100010011000;
		12'b010000010010: colour_data = 24'b110010001100000011000000;
		12'b010000010011: colour_data = 24'b111010011110000111100001;
		12'b010000010100: colour_data = 24'b111010011110000111100001;
		12'b010000010101: colour_data = 24'b100001000111111101111111;

		12'b010000100000: colour_data = 24'b100001000111111101111111;
		12'b010000100001: colour_data = 24'b111010011110000111100001;
		12'b010000100010: colour_data = 24'b111010011110000111100001;
		12'b010000100011: colour_data = 24'b110010001100000011000000;
		12'b010000100100: colour_data = 24'b100111011001100010011000;
		12'b010000100101: colour_data = 24'b100111011001100010011000;
		12'b010000100110: colour_data = 24'b100111011001100010011000;
		12'b010000100111: colour_data = 24'b100111011001100010011000;
		12'b010000101000: colour_data = 24'b100111011001100010011000;
		12'b010000101001: colour_data = 24'b111010011110000111100001;
		12'b010000101010: colour_data = 24'b111010011110000111100001;
		12'b010000101011: colour_data = 24'b111010011110000111100001;
		12'b010000101100: colour_data = 24'b111010011110000111100001;
		12'b010000101101: colour_data = 24'b100111011001100010011000;
		12'b010000101110: colour_data = 24'b100111011001100010011000;
		12'b010000101111: colour_data = 24'b100111011001100010011000;
		12'b010000110000: colour_data = 24'b100111011001100010011000;
		12'b010000110001: colour_data = 24'b100111011001100010011000;
		12'b010000110010: colour_data = 24'b100111011001100010011000;
		12'b010000110011: colour_data = 24'b110010001100000011000000;
		12'b010000110100: colour_data = 24'b111010011110000111100001;
		12'b010000110101: colour_data = 24'b100001000111111101111111;

		12'b010001000000: colour_data = 24'b100001000111111101111111;
		12'b010001000001: colour_data = 24'b111010011110000111100001;
		12'b010001000010: colour_data = 24'b111010011110000111100001;
		12'b010001000011: colour_data = 24'b100111011001100010011000;
		12'b010001000100: colour_data = 24'b111010011110000111100001;
		12'b010001000101: colour_data = 24'b111111111111111111111111;
		12'b010001000110: colour_data = 24'b111111111111111111111111;
		12'b010001000111: colour_data = 24'b111111111111111111111111;
		12'b010001001000: colour_data = 24'b111010011110000111100001;
		12'b010001001001: colour_data = 24'b100111011001100010011000;
		12'b010001001010: colour_data = 24'b111010011110000111100001;
		12'b010001001011: colour_data = 24'b111010011110000111100001;
		12'b010001001100: colour_data = 24'b100111011001100010011000;
		12'b010001001101: colour_data = 24'b111010011110000111100001;
		12'b010001001110: colour_data = 24'b111010011110000111100001;
		12'b010001001111: colour_data = 24'b111010011110000111100001;
		12'b010001010000: colour_data = 24'b111010011110000111100001;
		12'b010001010001: colour_data = 24'b111010011110000111100001;
		12'b010001010010: colour_data = 24'b111010011110000111100001;
		12'b010001010011: colour_data = 24'b100111011001100010011000;
		12'b010001010100: colour_data = 24'b111010011110000111100001;
		12'b010001010101: colour_data = 24'b100001000111111101111111;

		12'b010001100000: colour_data = 24'b100001000111111101111111;
		12'b010001100001: colour_data = 24'b110010001100000011000000;
		12'b010001100010: colour_data = 24'b111010011110000111100001;
		12'b010001100011: colour_data = 24'b100111011001100010011000;
		12'b010001100100: colour_data = 24'b111111111111111111111111;
		12'b010001100101: colour_data = 24'b111111111111111111111111;
		12'b010001100110: colour_data = 24'b111111111111111111111111;
		12'b010001100111: colour_data = 24'b111111111111111111111111;
		12'b010001101000: colour_data = 24'b100111011001100010011000;
		12'b010001101001: colour_data = 24'b110010001100000011000000;
		12'b010001101010: colour_data = 24'b110010001100000011000000;
		12'b010001101011: colour_data = 24'b100111011001100010011000;
		12'b010001101100: colour_data = 24'b111010011110000111100001;
		12'b010001101101: colour_data = 24'b100111011001100010011000;
		12'b010001101110: colour_data = 24'b100111011001100010011000;
		12'b010001101111: colour_data = 24'b100111011001100010011000;
		12'b010001110000: colour_data = 24'b100111011001100010011000;
		12'b010001110001: colour_data = 24'b100111011001100010011000;
		12'b010001110010: colour_data = 24'b100111011001100010011000;
		12'b010001110011: colour_data = 24'b111111111111111111111111;
		12'b010001110100: colour_data = 24'b110010001100000011000000;
		12'b010001110101: colour_data = 24'b100001000111111101111111;

		12'b010010000000: colour_data = 24'b111111110000000010010110;
		12'b010010000001: colour_data = 24'b100001000111111101111111;
		12'b010010000010: colour_data = 24'b111010011110000111100001;
		12'b010010000011: colour_data = 24'b100111011001100010011000;
		12'b010010000100: colour_data = 24'b111111111111111111111111;
		12'b010010000101: colour_data = 24'b111111111111111111111111;
		12'b010010000110: colour_data = 24'b111010011110000111100001;
		12'b010010000111: colour_data = 24'b100111011001100010011000;
		12'b010010001000: colour_data = 24'b110010001100000011000000;
		12'b010010001001: colour_data = 24'b110010001100000011000000;
		12'b010010001010: colour_data = 24'b110010001100000011000000;
		12'b010010001011: colour_data = 24'b110010001100000011000000;
		12'b010010001100: colour_data = 24'b100111011001100010011000;
		12'b010010001101: colour_data = 24'b111010011110000111100001;
		12'b010010001110: colour_data = 24'b111010011110000111100001;
		12'b010010001111: colour_data = 24'b111010011110000111100001;
		12'b010010010000: colour_data = 24'b111010011110000111100001;
		12'b010010010001: colour_data = 24'b111010011110000111100001;
		12'b010010010010: colour_data = 24'b100111011001100010011000;
		12'b010010010011: colour_data = 24'b111010011110000111100001;
		12'b010010010100: colour_data = 24'b100001000111111101111111;
		12'b010010010101: colour_data = 24'b111111110000000010010110;

		12'b010010100000: colour_data = 24'b111111110000000010010110;
		12'b010010100001: colour_data = 24'b100001000111111101111111;
		12'b010010100010: colour_data = 24'b110010001100000011000000;
		12'b010010100011: colour_data = 24'b111111111111111111111111;
		12'b010010100100: colour_data = 24'b100111011001100010011000;
		12'b010010100101: colour_data = 24'b100111011001100010011000;
		12'b010010100110: colour_data = 24'b100111011001100010011000;
		12'b010010100111: colour_data = 24'b100111011001100010011000;
		12'b010010101000: colour_data = 24'b110010001100000011000000;
		12'b010010101001: colour_data = 24'b110010001100000011000000;
		12'b010010101010: colour_data = 24'b110010001100000011000000;
		12'b010010101011: colour_data = 24'b110010001100000011000000;
		12'b010010101100: colour_data = 24'b110010001100000011000000;
		12'b010010101101: colour_data = 24'b100111011001100010011000;
		12'b010010101110: colour_data = 24'b100111011001100010011000;
		12'b010010101111: colour_data = 24'b100111011001100010011000;
		12'b010010110000: colour_data = 24'b100111011001100010011000;
		12'b010010110001: colour_data = 24'b100111011001100010011000;
		12'b010010110010: colour_data = 24'b111111111111111111111111;
		12'b010010110011: colour_data = 24'b110010001100000011000000;
		12'b010010110100: colour_data = 24'b100001000111111101111111;
		12'b010010110101: colour_data = 24'b111111110000000010010110;

		12'b010011000000: colour_data = 24'b111111110000000010010110;
		12'b010011000001: colour_data = 24'b111111110000000010010110;
		12'b010011000010: colour_data = 24'b100001000111111101111111;
		12'b010011000011: colour_data = 24'b111010011110000111100001;
		12'b010011000100: colour_data = 24'b111111111111111111111111;
		12'b010011000101: colour_data = 24'b111111111111111111111111;
		12'b010011000110: colour_data = 24'b111111111111111111111111;
		12'b010011000111: colour_data = 24'b111111111111111111111111;
		12'b010011001000: colour_data = 24'b100111011001100010011000;
		12'b010011001001: colour_data = 24'b100111011001100010011000;
		12'b010011001010: colour_data = 24'b100111011001100010011000;
		12'b010011001011: colour_data = 24'b100111011001100010011000;
		12'b010011001100: colour_data = 24'b100111011001100010011000;
		12'b010011001101: colour_data = 24'b111111111111111111111111;
		12'b010011001110: colour_data = 24'b111111111111111111111111;
		12'b010011001111: colour_data = 24'b111111111111111111111111;
		12'b010011010000: colour_data = 24'b111111111111111111111111;
		12'b010011010001: colour_data = 24'b111111111111111111111111;
		12'b010011010010: colour_data = 24'b111010011110000111100001;
		12'b010011010011: colour_data = 24'b100001000111111101111111;
		12'b010011010100: colour_data = 24'b111111110000000010010110;
		12'b010011010101: colour_data = 24'b111111110000000010010110;

		12'b010011100000: colour_data = 24'b111111110000000010010110;
		12'b010011100001: colour_data = 24'b111111110000000010010110;
		12'b010011100010: colour_data = 24'b100001000111111101111111;
		12'b010011100011: colour_data = 24'b110010001100000011000000;
		12'b010011100100: colour_data = 24'b111010011110000111100001;
		12'b010011100101: colour_data = 24'b111010011110000111100001;
		12'b010011100110: colour_data = 24'b111010011110000111100001;
		12'b010011100111: colour_data = 24'b111010011110000111100001;
		12'b010011101000: colour_data = 24'b111111111111111111111111;
		12'b010011101001: colour_data = 24'b111111111111111111111111;
		12'b010011101010: colour_data = 24'b111111111111111111111111;
		12'b010011101011: colour_data = 24'b111111111111111111111111;
		12'b010011101100: colour_data = 24'b111111111111111111111111;
		12'b010011101101: colour_data = 24'b111010011110000111100001;
		12'b010011101110: colour_data = 24'b111010011110000111100001;
		12'b010011101111: colour_data = 24'b111010011110000111100001;
		12'b010011110000: colour_data = 24'b111010011110000111100001;
		12'b010011110001: colour_data = 24'b111010011110000111100001;
		12'b010011110010: colour_data = 24'b110010001100000011000000;
		12'b010011110011: colour_data = 24'b100001000111111101111111;
		12'b010011110100: colour_data = 24'b111111110000000010010110;
		12'b010011110101: colour_data = 24'b111111110000000010010110;

		12'b010100000000: colour_data = 24'b111111110000000010010110;
		12'b010100000001: colour_data = 24'b111111110000000010010110;
		12'b010100000010: colour_data = 24'b111111110000000010010110;
		12'b010100000011: colour_data = 24'b100001000111111101111111;
		12'b010100000100: colour_data = 24'b110010001100000011000000;
		12'b010100000101: colour_data = 24'b110010001100000011000000;
		12'b010100000110: colour_data = 24'b111010011110000111100001;
		12'b010100000111: colour_data = 24'b111010011110000111100001;
		12'b010100001000: colour_data = 24'b111010011110000111100001;
		12'b010100001001: colour_data = 24'b111010011110000111100001;
		12'b010100001010: colour_data = 24'b111010011110000111100001;
		12'b010100001011: colour_data = 24'b111010011110000111100001;
		12'b010100001100: colour_data = 24'b111010011110000111100001;
		12'b010100001101: colour_data = 24'b111010011110000111100001;
		12'b010100001110: colour_data = 24'b111010011110000111100001;
		12'b010100001111: colour_data = 24'b111010011110000111100001;
		12'b010100010000: colour_data = 24'b110010001100000011000000;
		12'b010100010001: colour_data = 24'b110010001100000011000000;
		12'b010100010010: colour_data = 24'b100001000111111101111111;
		12'b010100010011: colour_data = 24'b111111110000000010010110;
		12'b010100010100: colour_data = 24'b111111110000000010010110;
		12'b010100010101: colour_data = 24'b111111110000000010010110;

		12'b010100100000: colour_data = 24'b111111110000000010010110;
		12'b010100100001: colour_data = 24'b111111110000000010010110;
		12'b010100100010: colour_data = 24'b111111110000000010010110;
		12'b010100100011: colour_data = 24'b111111110000000010010110;
		12'b010100100100: colour_data = 24'b100001000111111101111111;
		12'b010100100101: colour_data = 24'b100001000111111101111111;
		12'b010100100110: colour_data = 24'b110010001100000011000000;
		12'b010100100111: colour_data = 24'b110010001100000011000000;
		12'b010100101000: colour_data = 24'b111010011110000111100001;
		12'b010100101001: colour_data = 24'b111010011110000111100001;
		12'b010100101010: colour_data = 24'b111010011110000111100001;
		12'b010100101011: colour_data = 24'b111010011110000111100001;
		12'b010100101100: colour_data = 24'b111010011110000111100001;
		12'b010100101101: colour_data = 24'b111010011110000111100001;
		12'b010100101110: colour_data = 24'b110010001100000011000000;
		12'b010100101111: colour_data = 24'b110010001100000011000000;
		12'b010100110000: colour_data = 24'b100001000111111101111111;
		12'b010100110001: colour_data = 24'b100001000111111101111111;
		12'b010100110010: colour_data = 24'b111111110000000010010110;
		12'b010100110011: colour_data = 24'b111111110000000010010110;
		12'b010100110100: colour_data = 24'b111111110000000010010110;
		12'b010100110101: colour_data = 24'b111111110000000010010110;

		12'b010101000000: colour_data = 24'b111111110000000010010110;
		12'b010101000001: colour_data = 24'b111111110000000010010110;
		12'b010101000010: colour_data = 24'b111111110000000010010110;
		12'b010101000011: colour_data = 24'b111111110000000010010110;
		12'b010101000100: colour_data = 24'b111111110000000010010110;
		12'b010101000101: colour_data = 24'b111111110000000010010110;
		12'b010101000110: colour_data = 24'b100001000111111101111111;
		12'b010101000111: colour_data = 24'b100001000111111101111111;
		12'b010101001000: colour_data = 24'b110010001100000011000000;
		12'b010101001001: colour_data = 24'b110010001100000011000000;
		12'b010101001010: colour_data = 24'b110010001100000011000000;
		12'b010101001011: colour_data = 24'b110010001100000011000000;
		12'b010101001100: colour_data = 24'b110010001100000011000000;
		12'b010101001101: colour_data = 24'b110010001100000011000000;
		12'b010101001110: colour_data = 24'b100001000111111101111111;
		12'b010101001111: colour_data = 24'b100001000111111101111111;
		12'b010101010000: colour_data = 24'b111111110000000010010110;
		12'b010101010001: colour_data = 24'b111111110000000010010110;
		12'b010101010010: colour_data = 24'b111111110000000010010110;
		12'b010101010011: colour_data = 24'b111111110000000010010110;
		12'b010101010100: colour_data = 24'b111111110000000010010110;
		12'b010101010101: colour_data = 24'b111111110000000010010110;

		12'b010101100000: colour_data = 24'b111111110000000010010110;
		12'b010101100001: colour_data = 24'b111111110000000010010110;
		12'b010101100010: colour_data = 24'b111111110000000010010110;
		12'b010101100011: colour_data = 24'b111111110000000010010110;
		12'b010101100100: colour_data = 24'b111111110000000010010110;
		12'b010101100101: colour_data = 24'b111111110000000010010110;
		12'b010101100110: colour_data = 24'b111111110000000010010110;
		12'b010101100111: colour_data = 24'b111111110000000010010110;
		12'b010101101000: colour_data = 24'b100001000111111101111111;
		12'b010101101001: colour_data = 24'b100001000111111101111111;
		12'b010101101010: colour_data = 24'b100001000111111101111111;
		12'b010101101011: colour_data = 24'b100001000111111101111111;
		12'b010101101100: colour_data = 24'b100001000111111101111111;
		12'b010101101101: colour_data = 24'b100001000111111101111111;
		12'b010101101110: colour_data = 24'b111111110000000010010110;
		12'b010101101111: colour_data = 24'b111111110000000010010110;
		12'b010101110000: colour_data = 24'b111111110000000010010110;
		12'b010101110001: colour_data = 24'b111111110000000010010110;
		12'b010101110010: colour_data = 24'b111111110000000010010110;
		12'b010101110011: colour_data = 24'b111111110000000010010110;
		12'b010101110100: colour_data = 24'b111111110000000010010110;
		12'b010101110101: colour_data = 24'b111111110000000010010110;

		12'b010110000000: colour_data = 24'b111111110000000010010110;
		12'b010110000001: colour_data = 24'b111111110000000010010110;
		12'b010110000010: colour_data = 24'b111111110000000010010110;
		12'b010110000011: colour_data = 24'b111111110000000010010110;
		12'b010110000100: colour_data = 24'b111111110000000010010110;
		12'b010110000101: colour_data = 24'b111111110000000010010110;
		12'b010110000110: colour_data = 24'b111111110000000010010110;
		12'b010110000111: colour_data = 24'b111111110000000010010110;
		12'b010110001000: colour_data = 24'b101110011000000100101111;
		12'b010110001001: colour_data = 24'b101110011000000100101111;
		12'b010110001010: colour_data = 24'b101110011000000100101111;
		12'b010110001011: colour_data = 24'b101110011000000100101111;
		12'b010110001100: colour_data = 24'b101110011000000100101111;
		12'b010110001101: colour_data = 24'b101110011000000100101111;
		12'b010110001110: colour_data = 24'b111111110000000010010110;
		12'b010110001111: colour_data = 24'b111111110000000010010110;
		12'b010110010000: colour_data = 24'b111111110000000010010110;
		12'b010110010001: colour_data = 24'b111111110000000010010110;
		12'b010110010010: colour_data = 24'b111111110000000010010110;
		12'b010110010011: colour_data = 24'b111111110000000010010110;
		12'b010110010100: colour_data = 24'b111111110000000010010110;
		12'b010110010101: colour_data = 24'b111111110000000010010110;

		12'b010110100000: colour_data = 24'b111111110000000010010110;
		12'b010110100001: colour_data = 24'b111111110000000010010110;
		12'b010110100010: colour_data = 24'b111111110000000010010110;
		12'b010110100011: colour_data = 24'b111111110000000010010110;
		12'b010110100100: colour_data = 24'b111111110000000010010110;
		12'b010110100101: colour_data = 24'b111111110000000010010110;
		12'b010110100110: colour_data = 24'b101110011000000100101111;
		12'b010110100111: colour_data = 24'b101110011000000100101111;
		12'b010110101000: colour_data = 24'b111111111101101101011111;
		12'b010110101001: colour_data = 24'b111111111101101101011111;
		12'b010110101010: colour_data = 24'b111111111101101101011111;
		12'b010110101011: colour_data = 24'b111111111101101101011111;
		12'b010110101100: colour_data = 24'b111111111101101101011111;
		12'b010110101101: colour_data = 24'b111111111101101101011111;
		12'b010110101110: colour_data = 24'b101110011000000100101111;
		12'b010110101111: colour_data = 24'b101110011000000100101111;
		12'b010110110000: colour_data = 24'b111111110000000010010110;
		12'b010110110001: colour_data = 24'b111111110000000010010110;
		12'b010110110010: colour_data = 24'b111111110000000010010110;
		12'b010110110011: colour_data = 24'b111111110000000010010110;
		12'b010110110100: colour_data = 24'b111111110000000010010110;
		12'b010110110101: colour_data = 24'b111111110000000010010110;

		12'b010111000000: colour_data = 24'b111111110000000010010110;
		12'b010111000001: colour_data = 24'b111111110000000010010110;
		12'b010111000010: colour_data = 24'b111111110000000010010110;
		12'b010111000011: colour_data = 24'b111111110000000010010110;
		12'b010111000100: colour_data = 24'b101110011000000100101111;
		12'b010111000101: colour_data = 24'b101110011000000100101111;
		12'b010111000110: colour_data = 24'b111111111101101101011111;
		12'b010111000111: colour_data = 24'b111111111101101101011111;
		12'b010111001000: colour_data = 24'b111111111011000101000001;
		12'b010111001001: colour_data = 24'b111111111011000101000001;
		12'b010111001010: colour_data = 24'b111111111011000101000001;
		12'b010111001011: colour_data = 24'b111111111011000101000001;
		12'b010111001100: colour_data = 24'b111111111011000101000001;
		12'b010111001101: colour_data = 24'b111111111011000101000001;
		12'b010111001110: colour_data = 24'b111111111101101101011111;
		12'b010111001111: colour_data = 24'b111111111101101101011111;
		12'b010111010000: colour_data = 24'b101110011000000100101111;
		12'b010111010001: colour_data = 24'b101110011000000100101111;
		12'b010111010010: colour_data = 24'b111111110000000010010110;
		12'b010111010011: colour_data = 24'b111111110000000010010110;
		12'b010111010100: colour_data = 24'b111111110000000010010110;
		12'b010111010101: colour_data = 24'b111111110000000010010110;

		12'b010111100000: colour_data = 24'b111111110000000010010110;
		12'b010111100001: colour_data = 24'b111111110000000010010110;
		12'b010111100010: colour_data = 24'b111111110000000010010110;
		12'b010111100011: colour_data = 24'b101110011000000100101111;
		12'b010111100100: colour_data = 24'b111111111101101101011111;
		12'b010111100101: colour_data = 24'b111111111101101101011111;
		12'b010111100110: colour_data = 24'b111111111011000101000001;
		12'b010111100111: colour_data = 24'b111111111011000101000001;
		12'b010111101000: colour_data = 24'b111111111011000101000001;
		12'b010111101001: colour_data = 24'b111111111011000101000001;
		12'b010111101010: colour_data = 24'b111111111011000101000001;
		12'b010111101011: colour_data = 24'b111111111011000101000001;
		12'b010111101100: colour_data = 24'b111111111011000101000001;
		12'b010111101101: colour_data = 24'b111111111011000101000001;
		12'b010111101110: colour_data = 24'b111111111011000101000001;
		12'b010111101111: colour_data = 24'b111111111011000101000001;
		12'b010111110000: colour_data = 24'b111111111101101101011111;
		12'b010111110001: colour_data = 24'b111111111101101101011111;
		12'b010111110010: colour_data = 24'b101110011000000100101111;
		12'b010111110011: colour_data = 24'b111111110000000010010110;
		12'b010111110100: colour_data = 24'b111111110000000010010110;
		12'b010111110101: colour_data = 24'b111111110000000010010110;

		12'b011000000000: colour_data = 24'b111111110000000010010110;
		12'b011000000001: colour_data = 24'b111111110000000010010110;
		12'b011000000010: colour_data = 24'b101110011000000100101111;
		12'b011000000011: colour_data = 24'b111111111101101101011111;
		12'b011000000100: colour_data = 24'b111111111011000101000001;
		12'b011000000101: colour_data = 24'b111111111011000101000001;
		12'b011000000110: colour_data = 24'b111111111011000101000001;
		12'b011000000111: colour_data = 24'b111111111011000101000001;
		12'b011000001000: colour_data = 24'b111111111011000101000001;
		12'b011000001001: colour_data = 24'b111010101010001000111100;
		12'b011000001010: colour_data = 24'b111010101010001000111100;
		12'b011000001011: colour_data = 24'b111010101010001000111100;
		12'b011000001100: colour_data = 24'b111010101010001000111100;
		12'b011000001101: colour_data = 24'b111010101010001000111100;
		12'b011000001110: colour_data = 24'b111010101010001000111100;
		12'b011000001111: colour_data = 24'b111111111011000101000001;
		12'b011000010000: colour_data = 24'b111111111011000101000001;
		12'b011000010001: colour_data = 24'b111111111011000101000001;
		12'b011000010010: colour_data = 24'b111111111101101101011111;
		12'b011000010011: colour_data = 24'b101110011000000100101111;
		12'b011000010100: colour_data = 24'b111111110000000010010110;
		12'b011000010101: colour_data = 24'b111111110000000010010110;

		12'b011000100000: colour_data = 24'b111111110000000010010110;
		12'b011000100001: colour_data = 24'b111111110000000010010110;
		12'b011000100010: colour_data = 24'b101110011000000100101111;
		12'b011000100011: colour_data = 24'b111111111011000101000001;
		12'b011000100100: colour_data = 24'b111111111011000101000001;
		12'b011000100101: colour_data = 24'b111111111011000101000001;
		12'b011000100110: colour_data = 24'b111111111011000101000001;
		12'b011000100111: colour_data = 24'b111010101010001000111100;
		12'b011000101000: colour_data = 24'b111010101010001000111100;
		12'b011000101001: colour_data = 24'b110110011001011100110111;
		12'b011000101010: colour_data = 24'b110110011001011100110111;
		12'b011000101011: colour_data = 24'b110110011001011100110111;
		12'b011000101100: colour_data = 24'b110110011001011100110111;
		12'b011000101101: colour_data = 24'b110110011001011100110111;
		12'b011000101110: colour_data = 24'b110110011001011100110111;
		12'b011000101111: colour_data = 24'b111010101010001000111100;
		12'b011000110000: colour_data = 24'b111111111011000101000001;
		12'b011000110001: colour_data = 24'b111111111011000101000001;
		12'b011000110010: colour_data = 24'b111111111011000101000001;
		12'b011000110011: colour_data = 24'b101110011000000100101111;
		12'b011000110100: colour_data = 24'b111111110000000010010110;
		12'b011000110101: colour_data = 24'b111111110000000010010110;

		12'b011001000000: colour_data = 24'b111111110000000010010110;
		12'b011001000001: colour_data = 24'b101110011000000100101111;
		12'b011001000010: colour_data = 24'b111111111101101101011111;
		12'b011001000011: colour_data = 24'b111111111011000101000001;
		12'b011001000100: colour_data = 24'b111111111011000101000001;
		12'b011001000101: colour_data = 24'b111111111011000101000001;
		12'b011001000110: colour_data = 24'b111010101010001000111100;
		12'b011001000111: colour_data = 24'b110110011001011100110111;
		12'b011001001000: colour_data = 24'b110110011001011100110111;
		12'b011001001001: colour_data = 24'b111111111101101101011111;
		12'b011001001010: colour_data = 24'b111111111101101101011111;
		12'b011001001011: colour_data = 24'b111111111101101101011111;
		12'b011001001100: colour_data = 24'b110110011001011100110111;
		12'b011001001101: colour_data = 24'b111111111011000101000001;
		12'b011001001110: colour_data = 24'b111111111011000101000001;
		12'b011001001111: colour_data = 24'b110110011001011100110111;
		12'b011001010000: colour_data = 24'b111010101010001000111100;
		12'b011001010001: colour_data = 24'b111111111011000101000001;
		12'b011001010010: colour_data = 24'b111111111011000101000001;
		12'b011001010011: colour_data = 24'b111111111101101101011111;
		12'b011001010100: colour_data = 24'b101110011000000100101111;
		12'b011001010101: colour_data = 24'b111111110000000010010110;

		12'b011001100000: colour_data = 24'b111111110000000010010110;
		12'b011001100001: colour_data = 24'b101110011000000100101111;
		12'b011001100010: colour_data = 24'b111111111011000101000001;
		12'b011001100011: colour_data = 24'b111111111011000101000001;
		12'b011001100100: colour_data = 24'b111111111011000101000001;
		12'b011001100101: colour_data = 24'b111010101010001000111100;
		12'b011001100110: colour_data = 24'b110110011001011100110111;
		12'b011001100111: colour_data = 24'b111111111101101101011111;
		12'b011001101000: colour_data = 24'b111111111101101101011111;
		12'b011001101001: colour_data = 24'b111111111011000101000001;
		12'b011001101010: colour_data = 24'b111111111011000101000001;
		12'b011001101011: colour_data = 24'b110110011001011100110111;
		12'b011001101100: colour_data = 24'b111111111011000101000001;
		12'b011001101101: colour_data = 24'b111111111011000101000001;
		12'b011001101110: colour_data = 24'b111111111011000101000001;
		12'b011001101111: colour_data = 24'b111111111011000101000001;
		12'b011001110000: colour_data = 24'b110110011001011100110111;
		12'b011001110001: colour_data = 24'b111010101010001000111100;
		12'b011001110010: colour_data = 24'b111111111011000101000001;
		12'b011001110011: colour_data = 24'b111111111011000101000001;
		12'b011001110100: colour_data = 24'b101110011000000100101111;
		12'b011001110101: colour_data = 24'b111111110000000010010110;

		12'b011010000000: colour_data = 24'b101110011000000100101111;
		12'b011010000001: colour_data = 24'b111111111101101101011111;
		12'b011010000010: colour_data = 24'b111111111011000101000001;
		12'b011010000011: colour_data = 24'b111111111011000101000001;
		12'b011010000100: colour_data = 24'b111111111011000101000001;
		12'b011010000101: colour_data = 24'b110110011001011100110111;
		12'b011010000110: colour_data = 24'b111111111101101101011111;
		12'b011010000111: colour_data = 24'b111111111011000101000001;
		12'b011010001000: colour_data = 24'b111111111011000101000001;
		12'b011010001001: colour_data = 24'b111111111011000101000001;
		12'b011010001010: colour_data = 24'b111111111011000101000001;
		12'b011010001011: colour_data = 24'b110110011001011100110111;
		12'b011010001100: colour_data = 24'b111010101010001000111100;
		12'b011010001101: colour_data = 24'b111111111011000101000001;
		12'b011010001110: colour_data = 24'b111111111011000101000001;
		12'b011010001111: colour_data = 24'b110110011001011100110111;
		12'b011010010000: colour_data = 24'b111111111011000101000001;
		12'b011010010001: colour_data = 24'b110110011001011100110111;
		12'b011010010010: colour_data = 24'b111111111011000101000001;
		12'b011010010011: colour_data = 24'b111111111011000101000001;
		12'b011010010100: colour_data = 24'b111111111101101101011111;
		12'b011010010101: colour_data = 24'b101110011000000100101111;

		12'b011010100000: colour_data = 24'b101110011000000100101111;
		12'b011010100001: colour_data = 24'b111111111011000101000001;
		12'b011010100010: colour_data = 24'b111111111011000101000001;
		12'b011010100011: colour_data = 24'b111111111011000101000001;
		12'b011010100100: colour_data = 24'b110110011001011100110111;
		12'b011010100101: colour_data = 24'b111111111101101101011111;
		12'b011010100110: colour_data = 24'b111111111011000101000001;
		12'b011010100111: colour_data = 24'b111111111011000101000001;
		12'b011010101000: colour_data = 24'b111111111011000101000001;
		12'b011010101001: colour_data = 24'b111111111011000101000001;
		12'b011010101010: colour_data = 24'b111111111011000101000001;
		12'b011010101011: colour_data = 24'b110110011001011100110111;
		12'b011010101100: colour_data = 24'b111010101010001000111100;
		12'b011010101101: colour_data = 24'b111111111011000101000001;
		12'b011010101110: colour_data = 24'b111111111011000101000001;
		12'b011010101111: colour_data = 24'b110110011001011100110111;
		12'b011010110000: colour_data = 24'b111111111011000101000001;
		12'b011010110001: colour_data = 24'b110110011001011100110111;
		12'b011010110010: colour_data = 24'b111111111011000101000001;
		12'b011010110011: colour_data = 24'b111111111011000101000001;
		12'b011010110100: colour_data = 24'b111111111011000101000001;
		12'b011010110101: colour_data = 24'b101110011000000100101111;

		12'b011011000000: colour_data = 24'b101110011000000100101111;
		12'b011011000001: colour_data = 24'b111111111011000101000001;
		12'b011011000010: colour_data = 24'b111111111011000101000001;
		12'b011011000011: colour_data = 24'b111111111011000101000001;
		12'b011011000100: colour_data = 24'b110110011001011100110111;
		12'b011011000101: colour_data = 24'b111111111011000101000001;
		12'b011011000110: colour_data = 24'b111111111011000101000001;
		12'b011011000111: colour_data = 24'b111111111011000101000001;
		12'b011011001000: colour_data = 24'b111111111011000101000001;
		12'b011011001001: colour_data = 24'b111111111011000101000001;
		12'b011011001010: colour_data = 24'b111111111011000101000001;
		12'b011011001011: colour_data = 24'b111111111011000101000001;
		12'b011011001100: colour_data = 24'b110110011001011100110111;
		12'b011011001101: colour_data = 24'b111010101010001000111100;
		12'b011011001110: colour_data = 24'b111111111011000101000001;
		12'b011011001111: colour_data = 24'b111111111011000101000001;
		12'b011011010000: colour_data = 24'b111111111011000101000001;
		12'b011011010001: colour_data = 24'b110110011001011100110111;
		12'b011011010010: colour_data = 24'b111010101010001000111100;
		12'b011011010011: colour_data = 24'b111111111011000101000001;
		12'b011011010100: colour_data = 24'b111111111011000101000001;
		12'b011011010101: colour_data = 24'b101110011000000100101111;

		12'b011011100000: colour_data = 24'b101110011000000100101111;
		12'b011011100001: colour_data = 24'b111111111011000101000001;
		12'b011011100010: colour_data = 24'b111111111011000101000001;
		12'b011011100011: colour_data = 24'b111010101010001000111100;
		12'b011011100100: colour_data = 24'b110110011001011100110111;
		12'b011011100101: colour_data = 24'b110110011001011100110111;
		12'b011011100110: colour_data = 24'b110110011001011100110111;
		12'b011011100111: colour_data = 24'b110110011001011100110111;
		12'b011011101000: colour_data = 24'b110110011001011100110111;
		12'b011011101001: colour_data = 24'b111111111011000101000001;
		12'b011011101010: colour_data = 24'b111111111011000101000001;
		12'b011011101011: colour_data = 24'b111111111011000101000001;
		12'b011011101100: colour_data = 24'b111111111011000101000001;
		12'b011011101101: colour_data = 24'b110110011001011100110111;
		12'b011011101110: colour_data = 24'b110110011001011100110111;
		12'b011011101111: colour_data = 24'b110110011001011100110111;
		12'b011011110000: colour_data = 24'b110110011001011100110111;
		12'b011011110001: colour_data = 24'b110110011001011100110111;
		12'b011011110010: colour_data = 24'b110110011001011100110111;
		12'b011011110011: colour_data = 24'b111010101010001000111100;
		12'b011011110100: colour_data = 24'b111111111011000101000001;
		12'b011011110101: colour_data = 24'b101110011000000100101111;

		12'b011100000000: colour_data = 24'b101110011000000100101111;
		12'b011100000001: colour_data = 24'b111111111011000101000001;
		12'b011100000010: colour_data = 24'b111111111011000101000001;
		12'b011100000011: colour_data = 24'b110110011001011100110111;
		12'b011100000100: colour_data = 24'b111111111011000101000001;
		12'b011100000101: colour_data = 24'b111111111101101101011111;
		12'b011100000110: colour_data = 24'b111111111101101101011111;
		12'b011100000111: colour_data = 24'b111111111101101101011111;
		12'b011100001000: colour_data = 24'b111111111011000101000001;
		12'b011100001001: colour_data = 24'b110110011001011100110111;
		12'b011100001010: colour_data = 24'b111111111011000101000001;
		12'b011100001011: colour_data = 24'b111111111011000101000001;
		12'b011100001100: colour_data = 24'b110110011001011100110111;
		12'b011100001101: colour_data = 24'b111111111011000101000001;
		12'b011100001110: colour_data = 24'b111111111011000101000001;
		12'b011100001111: colour_data = 24'b111111111011000101000001;
		12'b011100010000: colour_data = 24'b111111111011000101000001;
		12'b011100010001: colour_data = 24'b111111111011000101000001;
		12'b011100010010: colour_data = 24'b111111111011000101000001;
		12'b011100010011: colour_data = 24'b110110011001011100110111;
		12'b011100010100: colour_data = 24'b111111111011000101000001;
		12'b011100010101: colour_data = 24'b101110011000000100101111;

		12'b011100100000: colour_data = 24'b101110011000000100101111;
		12'b011100100001: colour_data = 24'b111010101010001000111100;
		12'b011100100010: colour_data = 24'b111111111011000101000001;
		12'b011100100011: colour_data = 24'b110110011001011100110111;
		12'b011100100100: colour_data = 24'b111111111101101101011111;
		12'b011100100101: colour_data = 24'b111111111101101101011111;
		12'b011100100110: colour_data = 24'b111111111101101101011111;
		12'b011100100111: colour_data = 24'b111111111101101101011111;
		12'b011100101000: colour_data = 24'b110110011001011100110111;
		12'b011100101001: colour_data = 24'b111010101010001000111100;
		12'b011100101010: colour_data = 24'b111010101010001000111100;
		12'b011100101011: colour_data = 24'b110110011001011100110111;
		12'b011100101100: colour_data = 24'b111111111011000101000001;
		12'b011100101101: colour_data = 24'b110110011001011100110111;
		12'b011100101110: colour_data = 24'b110110011001011100110111;
		12'b011100101111: colour_data = 24'b110110011001011100110111;
		12'b011100110000: colour_data = 24'b110110011001011100110111;
		12'b011100110001: colour_data = 24'b110110011001011100110111;
		12'b011100110010: colour_data = 24'b110110011001011100110111;
		12'b011100110011: colour_data = 24'b111111111101101101011111;
		12'b011100110100: colour_data = 24'b111010101010001000111100;
		12'b011100110101: colour_data = 24'b101110011000000100101111;

		12'b011101000000: colour_data = 24'b111111110000000010010110;
		12'b011101000001: colour_data = 24'b101110011000000100101111;
		12'b011101000010: colour_data = 24'b111111111011000101000001;
		12'b011101000011: colour_data = 24'b110110011001011100110111;
		12'b011101000100: colour_data = 24'b111111111101101101011111;
		12'b011101000101: colour_data = 24'b111111111101101101011111;
		12'b011101000110: colour_data = 24'b111111111011000101000001;
		12'b011101000111: colour_data = 24'b110110011001011100110111;
		12'b011101001000: colour_data = 24'b111010101010001000111100;
		12'b011101001001: colour_data = 24'b111010101010001000111100;
		12'b011101001010: colour_data = 24'b111010101010001000111100;
		12'b011101001011: colour_data = 24'b111010101010001000111100;
		12'b011101001100: colour_data = 24'b110110011001011100110111;
		12'b011101001101: colour_data = 24'b111111111011000101000001;
		12'b011101001110: colour_data = 24'b111111111011000101000001;
		12'b011101001111: colour_data = 24'b111111111011000101000001;
		12'b011101010000: colour_data = 24'b111111111011000101000001;
		12'b011101010001: colour_data = 24'b111111111011000101000001;
		12'b011101010010: colour_data = 24'b110110011001011100110111;
		12'b011101010011: colour_data = 24'b111111111011000101000001;
		12'b011101010100: colour_data = 24'b101110011000000100101111;
		12'b011101010101: colour_data = 24'b111111110000000010010110;

		12'b011101100000: colour_data = 24'b111111110000000010010110;
		12'b011101100001: colour_data = 24'b101110011000000100101111;
		12'b011101100010: colour_data = 24'b111010101010001000111100;
		12'b011101100011: colour_data = 24'b111111111101101101011111;
		12'b011101100100: colour_data = 24'b110110011001011100110111;
		12'b011101100101: colour_data = 24'b110110011001011100110111;
		12'b011101100110: colour_data = 24'b110110011001011100110111;
		12'b011101100111: colour_data = 24'b110110011001011100110111;
		12'b011101101000: colour_data = 24'b111010101010001000111100;
		12'b011101101001: colour_data = 24'b111010101010001000111100;
		12'b011101101010: colour_data = 24'b111010101010001000111100;
		12'b011101101011: colour_data = 24'b111010101010001000111100;
		12'b011101101100: colour_data = 24'b111010101010001000111100;
		12'b011101101101: colour_data = 24'b110110011001011100110111;
		12'b011101101110: colour_data = 24'b110110011001011100110111;
		12'b011101101111: colour_data = 24'b110110011001011100110111;
		12'b011101110000: colour_data = 24'b110110011001011100110111;
		12'b011101110001: colour_data = 24'b110110011001011100110111;
		12'b011101110010: colour_data = 24'b111111111101101101011111;
		12'b011101110011: colour_data = 24'b111010101010001000111100;
		12'b011101110100: colour_data = 24'b101110011000000100101111;
		12'b011101110101: colour_data = 24'b111111110000000010010110;

		12'b011110000000: colour_data = 24'b111111110000000010010110;
		12'b011110000001: colour_data = 24'b111111110000000010010110;
		12'b011110000010: colour_data = 24'b101110011000000100101111;
		12'b011110000011: colour_data = 24'b111111111011000101000001;
		12'b011110000100: colour_data = 24'b111111111101101101011111;
		12'b011110000101: colour_data = 24'b111111111101101101011111;
		12'b011110000110: colour_data = 24'b111111111101101101011111;
		12'b011110000111: colour_data = 24'b111111111101101101011111;
		12'b011110001000: colour_data = 24'b110110011001011100110111;
		12'b011110001001: colour_data = 24'b110110011001011100110111;
		12'b011110001010: colour_data = 24'b110110011001011100110111;
		12'b011110001011: colour_data = 24'b110110011001011100110111;
		12'b011110001100: colour_data = 24'b110110011001011100110111;
		12'b011110001101: colour_data = 24'b111111111101101101011111;
		12'b011110001110: colour_data = 24'b111111111101101101011111;
		12'b011110001111: colour_data = 24'b111111111101101101011111;
		12'b011110010000: colour_data = 24'b111111111101101101011111;
		12'b011110010001: colour_data = 24'b111111111101101101011111;
		12'b011110010010: colour_data = 24'b111111111011000101000001;
		12'b011110010011: colour_data = 24'b101110011000000100101111;
		12'b011110010100: colour_data = 24'b111111110000000010010110;
		12'b011110010101: colour_data = 24'b111111110000000010010110;

		12'b011110100000: colour_data = 24'b111111110000000010010110;
		12'b011110100001: colour_data = 24'b111111110000000010010110;
		12'b011110100010: colour_data = 24'b101110011000000100101111;
		12'b011110100011: colour_data = 24'b111010101010001000111100;
		12'b011110100100: colour_data = 24'b111111111011000101000001;
		12'b011110100101: colour_data = 24'b111111111011000101000001;
		12'b011110100110: colour_data = 24'b111111111011000101000001;
		12'b011110100111: colour_data = 24'b111111111011000101000001;
		12'b011110101000: colour_data = 24'b111111111101101101011111;
		12'b011110101001: colour_data = 24'b111111111101101101011111;
		12'b011110101010: colour_data = 24'b111111111101101101011111;
		12'b011110101011: colour_data = 24'b111111111101101101011111;
		12'b011110101100: colour_data = 24'b111111111101101101011111;
		12'b011110101101: colour_data = 24'b111111111011000101000001;
		12'b011110101110: colour_data = 24'b111111111011000101000001;
		12'b011110101111: colour_data = 24'b111111111011000101000001;
		12'b011110110000: colour_data = 24'b111111111011000101000001;
		12'b011110110001: colour_data = 24'b111111111011000101000001;
		12'b011110110010: colour_data = 24'b111010101010001000111100;
		12'b011110110011: colour_data = 24'b101110011000000100101111;
		12'b011110110100: colour_data = 24'b111111110000000010010110;
		12'b011110110101: colour_data = 24'b111111110000000010010110;

		12'b011111000000: colour_data = 24'b111111110000000010010110;
		12'b011111000001: colour_data = 24'b111111110000000010010110;
		12'b011111000010: colour_data = 24'b111111110000000010010110;
		12'b011111000011: colour_data = 24'b101110011000000100101111;
		12'b011111000100: colour_data = 24'b111010101010001000111100;
		12'b011111000101: colour_data = 24'b111010101010001000111100;
		12'b011111000110: colour_data = 24'b111111111011000101000001;
		12'b011111000111: colour_data = 24'b111111111011000101000001;
		12'b011111001000: colour_data = 24'b111111111011000101000001;
		12'b011111001001: colour_data = 24'b111111111011000101000001;
		12'b011111001010: colour_data = 24'b111111111011000101000001;
		12'b011111001011: colour_data = 24'b111111111011000101000001;
		12'b011111001100: colour_data = 24'b111111111011000101000001;
		12'b011111001101: colour_data = 24'b111111111011000101000001;
		12'b011111001110: colour_data = 24'b111111111011000101000001;
		12'b011111001111: colour_data = 24'b111111111011000101000001;
		12'b011111010000: colour_data = 24'b111010101010001000111100;
		12'b011111010001: colour_data = 24'b111010101010001000111100;
		12'b011111010010: colour_data = 24'b101110011000000100101111;
		12'b011111010011: colour_data = 24'b111111110000000010010110;
		12'b011111010100: colour_data = 24'b111111110000000010010110;
		12'b011111010101: colour_data = 24'b111111110000000010010110;

		12'b011111100000: colour_data = 24'b111111110000000010010110;
		12'b011111100001: colour_data = 24'b111111110000000010010110;
		12'b011111100010: colour_data = 24'b111111110000000010010110;
		12'b011111100011: colour_data = 24'b111111110000000010010110;
		12'b011111100100: colour_data = 24'b101110011000000100101111;
		12'b011111100101: colour_data = 24'b101110011000000100101111;
		12'b011111100110: colour_data = 24'b111010101010001000111100;
		12'b011111100111: colour_data = 24'b111010101010001000111100;
		12'b011111101000: colour_data = 24'b111111111011000101000001;
		12'b011111101001: colour_data = 24'b111111111011000101000001;
		12'b011111101010: colour_data = 24'b111111111011000101000001;
		12'b011111101011: colour_data = 24'b111111111011000101000001;
		12'b011111101100: colour_data = 24'b111111111011000101000001;
		12'b011111101101: colour_data = 24'b111111111011000101000001;
		12'b011111101110: colour_data = 24'b111010101010001000111100;
		12'b011111101111: colour_data = 24'b111010101010001000111100;
		12'b011111110000: colour_data = 24'b101110011000000100101111;
		12'b011111110001: colour_data = 24'b101110011000000100101111;
		12'b011111110010: colour_data = 24'b111111110000000010010110;
		12'b011111110011: colour_data = 24'b111111110000000010010110;
		12'b011111110100: colour_data = 24'b111111110000000010010110;
		12'b011111110101: colour_data = 24'b111111110000000010010110;

		12'b100000000000: colour_data = 24'b111111110000000010010110;
		12'b100000000001: colour_data = 24'b111111110000000010010110;
		12'b100000000010: colour_data = 24'b111111110000000010010110;
		12'b100000000011: colour_data = 24'b111111110000000010010110;
		12'b100000000100: colour_data = 24'b111111110000000010010110;
		12'b100000000101: colour_data = 24'b111111110000000010010110;
		12'b100000000110: colour_data = 24'b101110011000000100101111;
		12'b100000000111: colour_data = 24'b101110011000000100101111;
		12'b100000001000: colour_data = 24'b111010101010001000111100;
		12'b100000001001: colour_data = 24'b111010101010001000111100;
		12'b100000001010: colour_data = 24'b111010101010001000111100;
		12'b100000001011: colour_data = 24'b111010101010001000111100;
		12'b100000001100: colour_data = 24'b111010101010001000111100;
		12'b100000001101: colour_data = 24'b111010101010001000111100;
		12'b100000001110: colour_data = 24'b101110011000000100101111;
		12'b100000001111: colour_data = 24'b101110011000000100101111;
		12'b100000010000: colour_data = 24'b111111110000000010010110;
		12'b100000010001: colour_data = 24'b111111110000000010010110;
		12'b100000010010: colour_data = 24'b111111110000000010010110;
		12'b100000010011: colour_data = 24'b111111110000000010010110;
		12'b100000010100: colour_data = 24'b111111110000000010010110;
		12'b100000010101: colour_data = 24'b111111110000000010010110;

		12'b100000100000: colour_data = 24'b111111110000000010010110;
		12'b100000100001: colour_data = 24'b111111110000000010010110;
		12'b100000100010: colour_data = 24'b111111110000000010010110;
		12'b100000100011: colour_data = 24'b111111110000000010010110;
		12'b100000100100: colour_data = 24'b111111110000000010010110;
		12'b100000100101: colour_data = 24'b111111110000000010010110;
		12'b100000100110: colour_data = 24'b111111110000000010010110;
		12'b100000100111: colour_data = 24'b111111110000000010010110;
		12'b100000101000: colour_data = 24'b101110011000000100101111;
		12'b100000101001: colour_data = 24'b101110011000000100101111;
		12'b100000101010: colour_data = 24'b101110011000000100101111;
		12'b100000101011: colour_data = 24'b101110011000000100101111;
		12'b100000101100: colour_data = 24'b101110011000000100101111;
		12'b100000101101: colour_data = 24'b101110011000000100101111;
		12'b100000101110: colour_data = 24'b111111110000000010010110;
		12'b100000101111: colour_data = 24'b111111110000000010010110;
		12'b100000110000: colour_data = 24'b111111110000000010010110;
		12'b100000110001: colour_data = 24'b111111110000000010010110;
		12'b100000110010: colour_data = 24'b111111110000000010010110;
		12'b100000110011: colour_data = 24'b111111110000000010010110;
		12'b100000110100: colour_data = 24'b111111110000000010010110;
		12'b100000110101: colour_data = 24'b111111110000000010010110;

		default: colour_data = 24'b000000000000000000000000;
	endcase
endmodule